** sch_path: /foss/designs/sky130_op_amp/runs/RUN_2025-10-21_19-17-39/parameters/slew_rate/run_74/transient.sch
**.subckt transient
I0 VDD IBIAS 4.9999999999999996e-06
C1 Vout GND 2.5e-11 m=1
V0 VSS GND 0
V2 VDD GND 1.9
Evdrv1 VN GND Vout GND 1
V3 VP GND DC 0 PWL(0 0 100n 0 100.1n -200000.00000000003)
x1 VDD IBIAS VN VP Vout VDD VSS sky130_op_amp
**** begin user architecture code



.control


    * Step function applied at time 100ns, save transient data
    tran 10n 20u
    set wr_singlescale
    * Measure slew rates
    meas tran sr max deriv(v(Vout))/1e6

    * Write measured slew rates to file
    let sr_val = $&sr
    echo $&sr_val > /foss/designs/sky130_op_amp/runs/RUN_2025-10-21_19-17-39/parameters/slew_rate/run_74/transient_74.data
.endc




.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice ss

.include /foss/designs/sky130_op_amp/netlist/rcx/sky130_op_amp.spice

.temp 130

.option SEED=12345

* Flag unsafe operating conditions (exceeds models' specified limits)
.option warn=1


**** end user architecture code
**.ends
.GLOBAL GND
.end
