** sch_path: /foss/designs/sky130_op_amp/runs/RUN_2025-10-21_18-48-36/parameters/slew_rate/run_07/transient.sch
**.subckt transient
I0 VDD IBIAS 4.9999999999999996e-06
C1 Vout GND 2.5e-11 m=1
V0 VSS GND 0
V2 VDD GND CACE{vdd}
Evdrv1 VN GND Vout GND 1
V3 VP GND DC 0 PWL(0 0 100n 0 100.1n CACE{vdd})
x1 VDD IBIAS VN VP Vout VDD VSS sky130_op_amp
**** begin user architecture code



.control


    * Step function applied at time 100ns, save transient data
    tran 10n 20u
    set wr_singlescale
    * Measure slew rates
    meas tran sr_pos max deriv(v(Vout))
    meas tran sr_neg min deriv(v(Vout))

    * Write measured slew rates to file
    let sr_pos_val = $&sr_pos
    let sr_neg_val = $&sr_neg
    echo $&sr_pos_val $&sr_neg_val > /foss/designs/sky130_op_amp/runs/RUN_2025-10-21_18-48-36/parameters/slew_rate/run_07/transient_7.data
.endc




.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice ss

.include /foss/designs/sky130_op_amp/netlist/rcx/sky130_op_amp.spice

.temp 27

.option SEED=12345

* Flag unsafe operating conditions (exceeds models' specified limits)
.option warn=1


**** end user architecture code
**.ends
.GLOBAL GND
.end
