magic
tech sky130A
magscale 1 2
timestamp 1761058420
<< nwell >>
rect -1389 8753 493 10699
rect 6859 7763 8741 11017
<< pwell >>
rect 2943 9219 5322 10899
rect 2943 9049 3029 9219
rect 5236 9049 5322 9219
rect 2943 8797 5322 9049
rect 2943 8627 3029 8797
rect 5236 8627 5322 8797
rect 2943 8208 5322 8627
rect -2348 3788 1578 8150
rect 3482 3985 6376 7511
rect 9715 7338 10376 7787
rect 8218 3992 10080 7100
<< nmos >>
rect 3129 10499 3329 10699
rect 3387 10499 3587 10699
rect 3645 10499 3845 10699
rect 3903 10499 4103 10699
rect 4161 10499 4361 10699
rect 4419 10499 4619 10699
rect 4677 10499 4877 10699
rect 4935 10499 5135 10699
rect 3129 10081 3329 10281
rect 3387 10081 3587 10281
rect 3645 10081 3845 10281
rect 3903 10081 4103 10281
rect 4161 10081 4361 10281
rect 4419 10081 4619 10281
rect 4677 10081 4877 10281
rect 4935 10081 5135 10281
rect 3129 9663 3329 9863
rect 3387 9663 3587 9863
rect 3645 9663 3845 9863
rect 3903 9663 4103 9863
rect 4161 9663 4361 9863
rect 4419 9663 4619 9863
rect 4677 9663 4877 9863
rect 4935 9663 5135 9863
rect 3129 9245 3329 9445
rect 3387 9245 3587 9445
rect 3645 9245 3845 9445
rect 3903 9245 4103 9445
rect 4161 9245 4361 9445
rect 4419 9245 4619 9445
rect 4677 9245 4877 9445
rect 4935 9245 5135 9445
rect 3129 8823 3329 9023
rect 3387 8823 3587 9023
rect 3645 8823 3845 9023
rect 3903 8823 4103 9023
rect 4161 8823 4361 9023
rect 4419 8823 4619 9023
rect 4677 8823 4877 9023
rect 4935 8823 5135 9023
rect 3129 8401 3329 8601
rect 3387 8401 3587 8601
rect 3645 8401 3845 8601
rect 3903 8401 4103 8601
rect 4161 8401 4361 8601
rect 4419 8401 4619 8601
rect 4677 8401 4877 8601
rect 4935 8401 5135 8601
rect -2162 7750 -1962 7950
rect -1904 7750 -1704 7950
rect -1646 7750 -1446 7950
rect -1388 7750 -1188 7950
rect -1130 7750 -930 7950
rect -872 7750 -672 7950
rect -614 7750 -414 7950
rect -356 7750 -156 7950
rect -98 7750 102 7950
rect 160 7750 360 7950
rect 418 7750 618 7950
rect 676 7750 876 7950
rect 934 7750 1134 7950
rect 1192 7750 1392 7950
rect -2162 7332 -1962 7532
rect -1904 7332 -1704 7532
rect -1646 7332 -1446 7532
rect -1388 7332 -1188 7532
rect -1130 7332 -930 7532
rect -872 7332 -672 7532
rect -614 7332 -414 7532
rect -356 7332 -156 7532
rect -98 7332 102 7532
rect 160 7332 360 7532
rect 418 7332 618 7532
rect 676 7332 876 7532
rect 934 7332 1134 7532
rect 1192 7332 1392 7532
rect -2162 6914 -1962 7114
rect -1904 6914 -1704 7114
rect -1646 6914 -1446 7114
rect -1388 6914 -1188 7114
rect -1130 6914 -930 7114
rect -872 6914 -672 7114
rect -614 6914 -414 7114
rect -356 6914 -156 7114
rect -98 6914 102 7114
rect 160 6914 360 7114
rect 418 6914 618 7114
rect 676 6914 876 7114
rect 934 6914 1134 7114
rect 1192 6914 1392 7114
rect -2162 6496 -1962 6696
rect -1904 6496 -1704 6696
rect -1646 6496 -1446 6696
rect -1388 6496 -1188 6696
rect -1130 6496 -930 6696
rect -872 6496 -672 6696
rect -614 6496 -414 6696
rect -356 6496 -156 6696
rect -98 6496 102 6696
rect 160 6496 360 6696
rect 418 6496 618 6696
rect 676 6496 876 6696
rect 934 6496 1134 6696
rect 1192 6496 1392 6696
rect -2162 6078 -1962 6278
rect -1904 6078 -1704 6278
rect -1646 6078 -1446 6278
rect -1388 6078 -1188 6278
rect -1130 6078 -930 6278
rect -872 6078 -672 6278
rect -614 6078 -414 6278
rect -356 6078 -156 6278
rect -98 6078 102 6278
rect 160 6078 360 6278
rect 418 6078 618 6278
rect 676 6078 876 6278
rect 934 6078 1134 6278
rect 1192 6078 1392 6278
rect -2162 5660 -1962 5860
rect -1904 5660 -1704 5860
rect -1646 5660 -1446 5860
rect -1388 5660 -1188 5860
rect -1130 5660 -930 5860
rect -872 5660 -672 5860
rect -614 5660 -414 5860
rect -356 5660 -156 5860
rect -98 5660 102 5860
rect 160 5660 360 5860
rect 418 5660 618 5860
rect 676 5660 876 5860
rect 934 5660 1134 5860
rect 1192 5660 1392 5860
rect -2162 5242 -1962 5442
rect -1904 5242 -1704 5442
rect -1646 5242 -1446 5442
rect -1388 5242 -1188 5442
rect -1130 5242 -930 5442
rect -872 5242 -672 5442
rect -614 5242 -414 5442
rect -356 5242 -156 5442
rect -98 5242 102 5442
rect 160 5242 360 5442
rect 418 5242 618 5442
rect 676 5242 876 5442
rect 934 5242 1134 5442
rect 1192 5242 1392 5442
rect -2162 4824 -1962 5024
rect -1904 4824 -1704 5024
rect -1646 4824 -1446 5024
rect -1388 4824 -1188 5024
rect -1130 4824 -930 5024
rect -872 4824 -672 5024
rect -614 4824 -414 5024
rect -356 4824 -156 5024
rect -98 4824 102 5024
rect 160 4824 360 5024
rect 418 4824 618 5024
rect 676 4824 876 5024
rect 934 4824 1134 5024
rect 1192 4824 1392 5024
rect -2162 4406 -1962 4606
rect -1904 4406 -1704 4606
rect -1646 4406 -1446 4606
rect -1388 4406 -1188 4606
rect -1130 4406 -930 4606
rect -872 4406 -672 4606
rect -614 4406 -414 4606
rect -356 4406 -156 4606
rect -98 4406 102 4606
rect 160 4406 360 4606
rect 418 4406 618 4606
rect 676 4406 876 4606
rect 934 4406 1134 4606
rect 1192 4406 1392 4606
rect -2162 3988 -1962 4188
rect -1904 3988 -1704 4188
rect -1646 3988 -1446 4188
rect -1388 3988 -1188 4188
rect -1130 3988 -930 4188
rect -872 3988 -672 4188
rect -614 3988 -414 4188
rect -356 3988 -156 4188
rect -98 3988 102 4188
rect 160 3988 360 4188
rect 418 3988 618 4188
rect 676 3988 876 4188
rect 934 3988 1134 4188
rect 1192 3988 1392 4188
rect 3668 7111 3868 7311
rect 3926 7111 4126 7311
rect 4184 7111 4384 7311
rect 4442 7111 4642 7311
rect 4700 7111 4900 7311
rect 4958 7111 5158 7311
rect 5216 7111 5416 7311
rect 5474 7111 5674 7311
rect 5732 7111 5932 7311
rect 5990 7111 6190 7311
rect 3668 6693 3868 6893
rect 3926 6693 4126 6893
rect 4184 6693 4384 6893
rect 4442 6693 4642 6893
rect 4700 6693 4900 6893
rect 4958 6693 5158 6893
rect 5216 6693 5416 6893
rect 5474 6693 5674 6893
rect 5732 6693 5932 6893
rect 5990 6693 6190 6893
rect 3668 6275 3868 6475
rect 3926 6275 4126 6475
rect 4184 6275 4384 6475
rect 4442 6275 4642 6475
rect 4700 6275 4900 6475
rect 4958 6275 5158 6475
rect 5216 6275 5416 6475
rect 5474 6275 5674 6475
rect 5732 6275 5932 6475
rect 5990 6275 6190 6475
rect 3668 5857 3868 6057
rect 3926 5857 4126 6057
rect 4184 5857 4384 6057
rect 4442 5857 4642 6057
rect 4700 5857 4900 6057
rect 4958 5857 5158 6057
rect 5216 5857 5416 6057
rect 5474 5857 5674 6057
rect 5732 5857 5932 6057
rect 5990 5857 6190 6057
rect 3668 5439 3868 5639
rect 3926 5439 4126 5639
rect 4184 5439 4384 5639
rect 4442 5439 4642 5639
rect 4700 5439 4900 5639
rect 4958 5439 5158 5639
rect 5216 5439 5416 5639
rect 5474 5439 5674 5639
rect 5732 5439 5932 5639
rect 5990 5439 6190 5639
rect 3668 5021 3868 5221
rect 3926 5021 4126 5221
rect 4184 5021 4384 5221
rect 4442 5021 4642 5221
rect 4700 5021 4900 5221
rect 4958 5021 5158 5221
rect 5216 5021 5416 5221
rect 5474 5021 5674 5221
rect 5732 5021 5932 5221
rect 5990 5021 6190 5221
rect 3668 4603 3868 4803
rect 3926 4603 4126 4803
rect 4184 4603 4384 4803
rect 4442 4603 4642 4803
rect 4700 4603 4900 4803
rect 4958 4603 5158 4803
rect 5216 4603 5416 4803
rect 5474 4603 5674 4803
rect 5732 4603 5932 4803
rect 5990 4603 6190 4803
rect 3668 4185 3868 4385
rect 3926 4185 4126 4385
rect 4184 4185 4384 4385
rect 4442 4185 4642 4385
rect 4700 4185 4900 4385
rect 4958 4185 5158 4385
rect 5216 4185 5416 4385
rect 5474 4185 5674 4385
rect 5732 4185 5932 4385
rect 5990 4185 6190 4385
rect 8404 6700 8604 6900
rect 8662 6700 8862 6900
rect 8920 6700 9120 6900
rect 9178 6700 9378 6900
rect 9436 6700 9636 6900
rect 9694 6700 9894 6900
rect 8404 6282 8604 6482
rect 8662 6282 8862 6482
rect 8920 6282 9120 6482
rect 9178 6282 9378 6482
rect 9436 6282 9636 6482
rect 9694 6282 9894 6482
rect 8404 5864 8604 6064
rect 8662 5864 8862 6064
rect 8920 5864 9120 6064
rect 9178 5864 9378 6064
rect 9436 5864 9636 6064
rect 9694 5864 9894 6064
rect 8404 5446 8604 5646
rect 8662 5446 8862 5646
rect 8920 5446 9120 5646
rect 9178 5446 9378 5646
rect 9436 5446 9636 5646
rect 9694 5446 9894 5646
rect 8404 5028 8604 5228
rect 8662 5028 8862 5228
rect 8920 5028 9120 5228
rect 9178 5028 9378 5228
rect 9436 5028 9636 5228
rect 9694 5028 9894 5228
rect 8404 4610 8604 4810
rect 8662 4610 8862 4810
rect 8920 4610 9120 4810
rect 9178 4610 9378 4810
rect 9436 4610 9636 4810
rect 9694 4610 9894 4810
rect 8404 4192 8604 4392
rect 8662 4192 8862 4392
rect 8920 4192 9120 4392
rect 9178 4192 9378 4392
rect 9436 4192 9636 4392
rect 9694 4192 9894 4392
<< pmos >>
rect -1193 10280 -993 10480
rect -935 10280 -735 10480
rect -677 10280 -477 10480
rect -419 10280 -219 10480
rect -161 10280 39 10480
rect 97 10280 297 10480
rect -1193 9844 -993 10044
rect -935 9844 -735 10044
rect -677 9844 -477 10044
rect -419 9844 -219 10044
rect -161 9844 39 10044
rect 97 9844 297 10044
rect -1193 9408 -993 9608
rect -935 9408 -735 9608
rect -677 9408 -477 9608
rect -419 9408 -219 9608
rect -161 9408 39 9608
rect 97 9408 297 9608
rect -1193 8972 -993 9172
rect -935 8972 -735 9172
rect -677 8972 -477 9172
rect -419 8972 -219 9172
rect -161 8972 39 9172
rect 97 8972 297 9172
rect 7055 10598 7255 10798
rect 7313 10598 7513 10798
rect 7571 10598 7771 10798
rect 7829 10598 8029 10798
rect 8087 10598 8287 10798
rect 8345 10598 8545 10798
rect 7055 10162 7255 10362
rect 7313 10162 7513 10362
rect 7571 10162 7771 10362
rect 7829 10162 8029 10362
rect 8087 10162 8287 10362
rect 8345 10162 8545 10362
rect 7055 9726 7255 9926
rect 7313 9726 7513 9926
rect 7571 9726 7771 9926
rect 7829 9726 8029 9926
rect 8087 9726 8287 9926
rect 8345 9726 8545 9926
rect 7055 9290 7255 9490
rect 7313 9290 7513 9490
rect 7571 9290 7771 9490
rect 7829 9290 8029 9490
rect 8087 9290 8287 9490
rect 8345 9290 8545 9490
rect 7055 8854 7255 9054
rect 7313 8854 7513 9054
rect 7571 8854 7771 9054
rect 7829 8854 8029 9054
rect 8087 8854 8287 9054
rect 8345 8854 8545 9054
rect 7055 8418 7255 8618
rect 7313 8418 7513 8618
rect 7571 8418 7771 8618
rect 7829 8418 8029 8618
rect 8087 8418 8287 8618
rect 8345 8418 8545 8618
rect 7055 7982 7255 8182
rect 7313 7982 7513 8182
rect 7571 7982 7771 8182
rect 7829 7982 8029 8182
rect 8087 7982 8287 8182
rect 8345 7982 8545 8182
<< ndiff >>
rect 3071 10684 3129 10699
rect 3071 10650 3083 10684
rect 3117 10650 3129 10684
rect 3071 10616 3129 10650
rect 3071 10582 3083 10616
rect 3117 10582 3129 10616
rect 3071 10548 3129 10582
rect 3071 10514 3083 10548
rect 3117 10514 3129 10548
rect 3071 10499 3129 10514
rect 3329 10684 3387 10699
rect 3329 10650 3341 10684
rect 3375 10650 3387 10684
rect 3329 10616 3387 10650
rect 3329 10582 3341 10616
rect 3375 10582 3387 10616
rect 3329 10548 3387 10582
rect 3329 10514 3341 10548
rect 3375 10514 3387 10548
rect 3329 10499 3387 10514
rect 3587 10684 3645 10699
rect 3587 10650 3599 10684
rect 3633 10650 3645 10684
rect 3587 10616 3645 10650
rect 3587 10582 3599 10616
rect 3633 10582 3645 10616
rect 3587 10548 3645 10582
rect 3587 10514 3599 10548
rect 3633 10514 3645 10548
rect 3587 10499 3645 10514
rect 3845 10684 3903 10699
rect 3845 10650 3857 10684
rect 3891 10650 3903 10684
rect 3845 10616 3903 10650
rect 3845 10582 3857 10616
rect 3891 10582 3903 10616
rect 3845 10548 3903 10582
rect 3845 10514 3857 10548
rect 3891 10514 3903 10548
rect 3845 10499 3903 10514
rect 4103 10684 4161 10699
rect 4103 10650 4115 10684
rect 4149 10650 4161 10684
rect 4103 10616 4161 10650
rect 4103 10582 4115 10616
rect 4149 10582 4161 10616
rect 4103 10548 4161 10582
rect 4103 10514 4115 10548
rect 4149 10514 4161 10548
rect 4103 10499 4161 10514
rect 4361 10684 4419 10699
rect 4361 10650 4373 10684
rect 4407 10650 4419 10684
rect 4361 10616 4419 10650
rect 4361 10582 4373 10616
rect 4407 10582 4419 10616
rect 4361 10548 4419 10582
rect 4361 10514 4373 10548
rect 4407 10514 4419 10548
rect 4361 10499 4419 10514
rect 4619 10684 4677 10699
rect 4619 10650 4631 10684
rect 4665 10650 4677 10684
rect 4619 10616 4677 10650
rect 4619 10582 4631 10616
rect 4665 10582 4677 10616
rect 4619 10548 4677 10582
rect 4619 10514 4631 10548
rect 4665 10514 4677 10548
rect 4619 10499 4677 10514
rect 4877 10684 4935 10699
rect 4877 10650 4889 10684
rect 4923 10650 4935 10684
rect 4877 10616 4935 10650
rect 4877 10582 4889 10616
rect 4923 10582 4935 10616
rect 4877 10548 4935 10582
rect 4877 10514 4889 10548
rect 4923 10514 4935 10548
rect 4877 10499 4935 10514
rect 5135 10684 5193 10699
rect 5135 10650 5147 10684
rect 5181 10650 5193 10684
rect 5135 10616 5193 10650
rect 5135 10582 5147 10616
rect 5181 10582 5193 10616
rect 5135 10548 5193 10582
rect 5135 10514 5147 10548
rect 5181 10514 5193 10548
rect 5135 10499 5193 10514
rect 3071 10266 3129 10281
rect 3071 10232 3083 10266
rect 3117 10232 3129 10266
rect 3071 10198 3129 10232
rect 3071 10164 3083 10198
rect 3117 10164 3129 10198
rect 3071 10130 3129 10164
rect 3071 10096 3083 10130
rect 3117 10096 3129 10130
rect 3071 10081 3129 10096
rect 3329 10266 3387 10281
rect 3329 10232 3341 10266
rect 3375 10232 3387 10266
rect 3329 10198 3387 10232
rect 3329 10164 3341 10198
rect 3375 10164 3387 10198
rect 3329 10130 3387 10164
rect 3329 10096 3341 10130
rect 3375 10096 3387 10130
rect 3329 10081 3387 10096
rect 3587 10266 3645 10281
rect 3587 10232 3599 10266
rect 3633 10232 3645 10266
rect 3587 10198 3645 10232
rect 3587 10164 3599 10198
rect 3633 10164 3645 10198
rect 3587 10130 3645 10164
rect 3587 10096 3599 10130
rect 3633 10096 3645 10130
rect 3587 10081 3645 10096
rect 3845 10266 3903 10281
rect 3845 10232 3857 10266
rect 3891 10232 3903 10266
rect 3845 10198 3903 10232
rect 3845 10164 3857 10198
rect 3891 10164 3903 10198
rect 3845 10130 3903 10164
rect 3845 10096 3857 10130
rect 3891 10096 3903 10130
rect 3845 10081 3903 10096
rect 4103 10266 4161 10281
rect 4103 10232 4115 10266
rect 4149 10232 4161 10266
rect 4103 10198 4161 10232
rect 4103 10164 4115 10198
rect 4149 10164 4161 10198
rect 4103 10130 4161 10164
rect 4103 10096 4115 10130
rect 4149 10096 4161 10130
rect 4103 10081 4161 10096
rect 4361 10266 4419 10281
rect 4361 10232 4373 10266
rect 4407 10232 4419 10266
rect 4361 10198 4419 10232
rect 4361 10164 4373 10198
rect 4407 10164 4419 10198
rect 4361 10130 4419 10164
rect 4361 10096 4373 10130
rect 4407 10096 4419 10130
rect 4361 10081 4419 10096
rect 4619 10266 4677 10281
rect 4619 10232 4631 10266
rect 4665 10232 4677 10266
rect 4619 10198 4677 10232
rect 4619 10164 4631 10198
rect 4665 10164 4677 10198
rect 4619 10130 4677 10164
rect 4619 10096 4631 10130
rect 4665 10096 4677 10130
rect 4619 10081 4677 10096
rect 4877 10266 4935 10281
rect 4877 10232 4889 10266
rect 4923 10232 4935 10266
rect 4877 10198 4935 10232
rect 4877 10164 4889 10198
rect 4923 10164 4935 10198
rect 4877 10130 4935 10164
rect 4877 10096 4889 10130
rect 4923 10096 4935 10130
rect 4877 10081 4935 10096
rect 5135 10266 5193 10281
rect 5135 10232 5147 10266
rect 5181 10232 5193 10266
rect 5135 10198 5193 10232
rect 5135 10164 5147 10198
rect 5181 10164 5193 10198
rect 5135 10130 5193 10164
rect 5135 10096 5147 10130
rect 5181 10096 5193 10130
rect 5135 10081 5193 10096
rect 3071 9848 3129 9863
rect 3071 9814 3083 9848
rect 3117 9814 3129 9848
rect 3071 9780 3129 9814
rect 3071 9746 3083 9780
rect 3117 9746 3129 9780
rect 3071 9712 3129 9746
rect 3071 9678 3083 9712
rect 3117 9678 3129 9712
rect 3071 9663 3129 9678
rect 3329 9848 3387 9863
rect 3329 9814 3341 9848
rect 3375 9814 3387 9848
rect 3329 9780 3387 9814
rect 3329 9746 3341 9780
rect 3375 9746 3387 9780
rect 3329 9712 3387 9746
rect 3329 9678 3341 9712
rect 3375 9678 3387 9712
rect 3329 9663 3387 9678
rect 3587 9848 3645 9863
rect 3587 9814 3599 9848
rect 3633 9814 3645 9848
rect 3587 9780 3645 9814
rect 3587 9746 3599 9780
rect 3633 9746 3645 9780
rect 3587 9712 3645 9746
rect 3587 9678 3599 9712
rect 3633 9678 3645 9712
rect 3587 9663 3645 9678
rect 3845 9848 3903 9863
rect 3845 9814 3857 9848
rect 3891 9814 3903 9848
rect 3845 9780 3903 9814
rect 3845 9746 3857 9780
rect 3891 9746 3903 9780
rect 3845 9712 3903 9746
rect 3845 9678 3857 9712
rect 3891 9678 3903 9712
rect 3845 9663 3903 9678
rect 4103 9848 4161 9863
rect 4103 9814 4115 9848
rect 4149 9814 4161 9848
rect 4103 9780 4161 9814
rect 4103 9746 4115 9780
rect 4149 9746 4161 9780
rect 4103 9712 4161 9746
rect 4103 9678 4115 9712
rect 4149 9678 4161 9712
rect 4103 9663 4161 9678
rect 4361 9848 4419 9863
rect 4361 9814 4373 9848
rect 4407 9814 4419 9848
rect 4361 9780 4419 9814
rect 4361 9746 4373 9780
rect 4407 9746 4419 9780
rect 4361 9712 4419 9746
rect 4361 9678 4373 9712
rect 4407 9678 4419 9712
rect 4361 9663 4419 9678
rect 4619 9848 4677 9863
rect 4619 9814 4631 9848
rect 4665 9814 4677 9848
rect 4619 9780 4677 9814
rect 4619 9746 4631 9780
rect 4665 9746 4677 9780
rect 4619 9712 4677 9746
rect 4619 9678 4631 9712
rect 4665 9678 4677 9712
rect 4619 9663 4677 9678
rect 4877 9848 4935 9863
rect 4877 9814 4889 9848
rect 4923 9814 4935 9848
rect 4877 9780 4935 9814
rect 4877 9746 4889 9780
rect 4923 9746 4935 9780
rect 4877 9712 4935 9746
rect 4877 9678 4889 9712
rect 4923 9678 4935 9712
rect 4877 9663 4935 9678
rect 5135 9848 5193 9863
rect 5135 9814 5147 9848
rect 5181 9814 5193 9848
rect 5135 9780 5193 9814
rect 5135 9746 5147 9780
rect 5181 9746 5193 9780
rect 5135 9712 5193 9746
rect 5135 9678 5147 9712
rect 5181 9678 5193 9712
rect 5135 9663 5193 9678
rect 3071 9430 3129 9445
rect 3071 9396 3083 9430
rect 3117 9396 3129 9430
rect 3071 9362 3129 9396
rect 3071 9328 3083 9362
rect 3117 9328 3129 9362
rect 3071 9294 3129 9328
rect 3071 9260 3083 9294
rect 3117 9260 3129 9294
rect 3071 9245 3129 9260
rect 3329 9430 3387 9445
rect 3329 9396 3341 9430
rect 3375 9396 3387 9430
rect 3329 9362 3387 9396
rect 3329 9328 3341 9362
rect 3375 9328 3387 9362
rect 3329 9294 3387 9328
rect 3329 9260 3341 9294
rect 3375 9260 3387 9294
rect 3329 9245 3387 9260
rect 3587 9430 3645 9445
rect 3587 9396 3599 9430
rect 3633 9396 3645 9430
rect 3587 9362 3645 9396
rect 3587 9328 3599 9362
rect 3633 9328 3645 9362
rect 3587 9294 3645 9328
rect 3587 9260 3599 9294
rect 3633 9260 3645 9294
rect 3587 9245 3645 9260
rect 3845 9430 3903 9445
rect 3845 9396 3857 9430
rect 3891 9396 3903 9430
rect 3845 9362 3903 9396
rect 3845 9328 3857 9362
rect 3891 9328 3903 9362
rect 3845 9294 3903 9328
rect 3845 9260 3857 9294
rect 3891 9260 3903 9294
rect 3845 9245 3903 9260
rect 4103 9430 4161 9445
rect 4103 9396 4115 9430
rect 4149 9396 4161 9430
rect 4103 9362 4161 9396
rect 4103 9328 4115 9362
rect 4149 9328 4161 9362
rect 4103 9294 4161 9328
rect 4103 9260 4115 9294
rect 4149 9260 4161 9294
rect 4103 9245 4161 9260
rect 4361 9430 4419 9445
rect 4361 9396 4373 9430
rect 4407 9396 4419 9430
rect 4361 9362 4419 9396
rect 4361 9328 4373 9362
rect 4407 9328 4419 9362
rect 4361 9294 4419 9328
rect 4361 9260 4373 9294
rect 4407 9260 4419 9294
rect 4361 9245 4419 9260
rect 4619 9430 4677 9445
rect 4619 9396 4631 9430
rect 4665 9396 4677 9430
rect 4619 9362 4677 9396
rect 4619 9328 4631 9362
rect 4665 9328 4677 9362
rect 4619 9294 4677 9328
rect 4619 9260 4631 9294
rect 4665 9260 4677 9294
rect 4619 9245 4677 9260
rect 4877 9430 4935 9445
rect 4877 9396 4889 9430
rect 4923 9396 4935 9430
rect 4877 9362 4935 9396
rect 4877 9328 4889 9362
rect 4923 9328 4935 9362
rect 4877 9294 4935 9328
rect 4877 9260 4889 9294
rect 4923 9260 4935 9294
rect 4877 9245 4935 9260
rect 5135 9430 5193 9445
rect 5135 9396 5147 9430
rect 5181 9396 5193 9430
rect 5135 9362 5193 9396
rect 5135 9328 5147 9362
rect 5181 9328 5193 9362
rect 5135 9294 5193 9328
rect 5135 9260 5147 9294
rect 5181 9260 5193 9294
rect 5135 9245 5193 9260
rect 3071 9008 3129 9023
rect 3071 8974 3083 9008
rect 3117 8974 3129 9008
rect 3071 8940 3129 8974
rect 3071 8906 3083 8940
rect 3117 8906 3129 8940
rect 3071 8872 3129 8906
rect 3071 8838 3083 8872
rect 3117 8838 3129 8872
rect 3071 8823 3129 8838
rect 3329 9008 3387 9023
rect 3329 8974 3341 9008
rect 3375 8974 3387 9008
rect 3329 8940 3387 8974
rect 3329 8906 3341 8940
rect 3375 8906 3387 8940
rect 3329 8872 3387 8906
rect 3329 8838 3341 8872
rect 3375 8838 3387 8872
rect 3329 8823 3387 8838
rect 3587 9008 3645 9023
rect 3587 8974 3599 9008
rect 3633 8974 3645 9008
rect 3587 8940 3645 8974
rect 3587 8906 3599 8940
rect 3633 8906 3645 8940
rect 3587 8872 3645 8906
rect 3587 8838 3599 8872
rect 3633 8838 3645 8872
rect 3587 8823 3645 8838
rect 3845 9008 3903 9023
rect 3845 8974 3857 9008
rect 3891 8974 3903 9008
rect 3845 8940 3903 8974
rect 3845 8906 3857 8940
rect 3891 8906 3903 8940
rect 3845 8872 3903 8906
rect 3845 8838 3857 8872
rect 3891 8838 3903 8872
rect 3845 8823 3903 8838
rect 4103 9008 4161 9023
rect 4103 8974 4115 9008
rect 4149 8974 4161 9008
rect 4103 8940 4161 8974
rect 4103 8906 4115 8940
rect 4149 8906 4161 8940
rect 4103 8872 4161 8906
rect 4103 8838 4115 8872
rect 4149 8838 4161 8872
rect 4103 8823 4161 8838
rect 4361 9008 4419 9023
rect 4361 8974 4373 9008
rect 4407 8974 4419 9008
rect 4361 8940 4419 8974
rect 4361 8906 4373 8940
rect 4407 8906 4419 8940
rect 4361 8872 4419 8906
rect 4361 8838 4373 8872
rect 4407 8838 4419 8872
rect 4361 8823 4419 8838
rect 4619 9008 4677 9023
rect 4619 8974 4631 9008
rect 4665 8974 4677 9008
rect 4619 8940 4677 8974
rect 4619 8906 4631 8940
rect 4665 8906 4677 8940
rect 4619 8872 4677 8906
rect 4619 8838 4631 8872
rect 4665 8838 4677 8872
rect 4619 8823 4677 8838
rect 4877 9008 4935 9023
rect 4877 8974 4889 9008
rect 4923 8974 4935 9008
rect 4877 8940 4935 8974
rect 4877 8906 4889 8940
rect 4923 8906 4935 8940
rect 4877 8872 4935 8906
rect 4877 8838 4889 8872
rect 4923 8838 4935 8872
rect 4877 8823 4935 8838
rect 5135 9008 5193 9023
rect 5135 8974 5147 9008
rect 5181 8974 5193 9008
rect 5135 8940 5193 8974
rect 5135 8906 5147 8940
rect 5181 8906 5193 8940
rect 5135 8872 5193 8906
rect 5135 8838 5147 8872
rect 5181 8838 5193 8872
rect 5135 8823 5193 8838
rect 3071 8586 3129 8601
rect 3071 8552 3083 8586
rect 3117 8552 3129 8586
rect 3071 8518 3129 8552
rect 3071 8484 3083 8518
rect 3117 8484 3129 8518
rect 3071 8450 3129 8484
rect 3071 8416 3083 8450
rect 3117 8416 3129 8450
rect 3071 8401 3129 8416
rect 3329 8586 3387 8601
rect 3329 8552 3341 8586
rect 3375 8552 3387 8586
rect 3329 8518 3387 8552
rect 3329 8484 3341 8518
rect 3375 8484 3387 8518
rect 3329 8450 3387 8484
rect 3329 8416 3341 8450
rect 3375 8416 3387 8450
rect 3329 8401 3387 8416
rect 3587 8586 3645 8601
rect 3587 8552 3599 8586
rect 3633 8552 3645 8586
rect 3587 8518 3645 8552
rect 3587 8484 3599 8518
rect 3633 8484 3645 8518
rect 3587 8450 3645 8484
rect 3587 8416 3599 8450
rect 3633 8416 3645 8450
rect 3587 8401 3645 8416
rect 3845 8586 3903 8601
rect 3845 8552 3857 8586
rect 3891 8552 3903 8586
rect 3845 8518 3903 8552
rect 3845 8484 3857 8518
rect 3891 8484 3903 8518
rect 3845 8450 3903 8484
rect 3845 8416 3857 8450
rect 3891 8416 3903 8450
rect 3845 8401 3903 8416
rect 4103 8586 4161 8601
rect 4103 8552 4115 8586
rect 4149 8552 4161 8586
rect 4103 8518 4161 8552
rect 4103 8484 4115 8518
rect 4149 8484 4161 8518
rect 4103 8450 4161 8484
rect 4103 8416 4115 8450
rect 4149 8416 4161 8450
rect 4103 8401 4161 8416
rect 4361 8586 4419 8601
rect 4361 8552 4373 8586
rect 4407 8552 4419 8586
rect 4361 8518 4419 8552
rect 4361 8484 4373 8518
rect 4407 8484 4419 8518
rect 4361 8450 4419 8484
rect 4361 8416 4373 8450
rect 4407 8416 4419 8450
rect 4361 8401 4419 8416
rect 4619 8586 4677 8601
rect 4619 8552 4631 8586
rect 4665 8552 4677 8586
rect 4619 8518 4677 8552
rect 4619 8484 4631 8518
rect 4665 8484 4677 8518
rect 4619 8450 4677 8484
rect 4619 8416 4631 8450
rect 4665 8416 4677 8450
rect 4619 8401 4677 8416
rect 4877 8586 4935 8601
rect 4877 8552 4889 8586
rect 4923 8552 4935 8586
rect 4877 8518 4935 8552
rect 4877 8484 4889 8518
rect 4923 8484 4935 8518
rect 4877 8450 4935 8484
rect 4877 8416 4889 8450
rect 4923 8416 4935 8450
rect 4877 8401 4935 8416
rect 5135 8586 5193 8601
rect 5135 8552 5147 8586
rect 5181 8552 5193 8586
rect 5135 8518 5193 8552
rect 5135 8484 5147 8518
rect 5181 8484 5193 8518
rect 5135 8450 5193 8484
rect 5135 8416 5147 8450
rect 5181 8416 5193 8450
rect 5135 8401 5193 8416
rect -2220 7935 -2162 7950
rect -2220 7901 -2208 7935
rect -2174 7901 -2162 7935
rect -2220 7867 -2162 7901
rect -2220 7833 -2208 7867
rect -2174 7833 -2162 7867
rect -2220 7799 -2162 7833
rect -2220 7765 -2208 7799
rect -2174 7765 -2162 7799
rect -2220 7750 -2162 7765
rect -1962 7935 -1904 7950
rect -1962 7901 -1950 7935
rect -1916 7901 -1904 7935
rect -1962 7867 -1904 7901
rect -1962 7833 -1950 7867
rect -1916 7833 -1904 7867
rect -1962 7799 -1904 7833
rect -1962 7765 -1950 7799
rect -1916 7765 -1904 7799
rect -1962 7750 -1904 7765
rect -1704 7935 -1646 7950
rect -1704 7901 -1692 7935
rect -1658 7901 -1646 7935
rect -1704 7867 -1646 7901
rect -1704 7833 -1692 7867
rect -1658 7833 -1646 7867
rect -1704 7799 -1646 7833
rect -1704 7765 -1692 7799
rect -1658 7765 -1646 7799
rect -1704 7750 -1646 7765
rect -1446 7935 -1388 7950
rect -1446 7901 -1434 7935
rect -1400 7901 -1388 7935
rect -1446 7867 -1388 7901
rect -1446 7833 -1434 7867
rect -1400 7833 -1388 7867
rect -1446 7799 -1388 7833
rect -1446 7765 -1434 7799
rect -1400 7765 -1388 7799
rect -1446 7750 -1388 7765
rect -1188 7935 -1130 7950
rect -1188 7901 -1176 7935
rect -1142 7901 -1130 7935
rect -1188 7867 -1130 7901
rect -1188 7833 -1176 7867
rect -1142 7833 -1130 7867
rect -1188 7799 -1130 7833
rect -1188 7765 -1176 7799
rect -1142 7765 -1130 7799
rect -1188 7750 -1130 7765
rect -930 7935 -872 7950
rect -930 7901 -918 7935
rect -884 7901 -872 7935
rect -930 7867 -872 7901
rect -930 7833 -918 7867
rect -884 7833 -872 7867
rect -930 7799 -872 7833
rect -930 7765 -918 7799
rect -884 7765 -872 7799
rect -930 7750 -872 7765
rect -672 7935 -614 7950
rect -672 7901 -660 7935
rect -626 7901 -614 7935
rect -672 7867 -614 7901
rect -672 7833 -660 7867
rect -626 7833 -614 7867
rect -672 7799 -614 7833
rect -672 7765 -660 7799
rect -626 7765 -614 7799
rect -672 7750 -614 7765
rect -414 7935 -356 7950
rect -414 7901 -402 7935
rect -368 7901 -356 7935
rect -414 7867 -356 7901
rect -414 7833 -402 7867
rect -368 7833 -356 7867
rect -414 7799 -356 7833
rect -414 7765 -402 7799
rect -368 7765 -356 7799
rect -414 7750 -356 7765
rect -156 7935 -98 7950
rect -156 7901 -144 7935
rect -110 7901 -98 7935
rect -156 7867 -98 7901
rect -156 7833 -144 7867
rect -110 7833 -98 7867
rect -156 7799 -98 7833
rect -156 7765 -144 7799
rect -110 7765 -98 7799
rect -156 7750 -98 7765
rect 102 7935 160 7950
rect 102 7901 114 7935
rect 148 7901 160 7935
rect 102 7867 160 7901
rect 102 7833 114 7867
rect 148 7833 160 7867
rect 102 7799 160 7833
rect 102 7765 114 7799
rect 148 7765 160 7799
rect 102 7750 160 7765
rect 360 7935 418 7950
rect 360 7901 372 7935
rect 406 7901 418 7935
rect 360 7867 418 7901
rect 360 7833 372 7867
rect 406 7833 418 7867
rect 360 7799 418 7833
rect 360 7765 372 7799
rect 406 7765 418 7799
rect 360 7750 418 7765
rect 618 7935 676 7950
rect 618 7901 630 7935
rect 664 7901 676 7935
rect 618 7867 676 7901
rect 618 7833 630 7867
rect 664 7833 676 7867
rect 618 7799 676 7833
rect 618 7765 630 7799
rect 664 7765 676 7799
rect 618 7750 676 7765
rect 876 7935 934 7950
rect 876 7901 888 7935
rect 922 7901 934 7935
rect 876 7867 934 7901
rect 876 7833 888 7867
rect 922 7833 934 7867
rect 876 7799 934 7833
rect 876 7765 888 7799
rect 922 7765 934 7799
rect 876 7750 934 7765
rect 1134 7935 1192 7950
rect 1134 7901 1146 7935
rect 1180 7901 1192 7935
rect 1134 7867 1192 7901
rect 1134 7833 1146 7867
rect 1180 7833 1192 7867
rect 1134 7799 1192 7833
rect 1134 7765 1146 7799
rect 1180 7765 1192 7799
rect 1134 7750 1192 7765
rect 1392 7935 1450 7950
rect 1392 7901 1404 7935
rect 1438 7901 1450 7935
rect 1392 7867 1450 7901
rect 1392 7833 1404 7867
rect 1438 7833 1450 7867
rect 1392 7799 1450 7833
rect 1392 7765 1404 7799
rect 1438 7765 1450 7799
rect 1392 7750 1450 7765
rect -2220 7517 -2162 7532
rect -2220 7483 -2208 7517
rect -2174 7483 -2162 7517
rect -2220 7449 -2162 7483
rect -2220 7415 -2208 7449
rect -2174 7415 -2162 7449
rect -2220 7381 -2162 7415
rect -2220 7347 -2208 7381
rect -2174 7347 -2162 7381
rect -2220 7332 -2162 7347
rect -1962 7517 -1904 7532
rect -1962 7483 -1950 7517
rect -1916 7483 -1904 7517
rect -1962 7449 -1904 7483
rect -1962 7415 -1950 7449
rect -1916 7415 -1904 7449
rect -1962 7381 -1904 7415
rect -1962 7347 -1950 7381
rect -1916 7347 -1904 7381
rect -1962 7332 -1904 7347
rect -1704 7517 -1646 7532
rect -1704 7483 -1692 7517
rect -1658 7483 -1646 7517
rect -1704 7449 -1646 7483
rect -1704 7415 -1692 7449
rect -1658 7415 -1646 7449
rect -1704 7381 -1646 7415
rect -1704 7347 -1692 7381
rect -1658 7347 -1646 7381
rect -1704 7332 -1646 7347
rect -1446 7517 -1388 7532
rect -1446 7483 -1434 7517
rect -1400 7483 -1388 7517
rect -1446 7449 -1388 7483
rect -1446 7415 -1434 7449
rect -1400 7415 -1388 7449
rect -1446 7381 -1388 7415
rect -1446 7347 -1434 7381
rect -1400 7347 -1388 7381
rect -1446 7332 -1388 7347
rect -1188 7517 -1130 7532
rect -1188 7483 -1176 7517
rect -1142 7483 -1130 7517
rect -1188 7449 -1130 7483
rect -1188 7415 -1176 7449
rect -1142 7415 -1130 7449
rect -1188 7381 -1130 7415
rect -1188 7347 -1176 7381
rect -1142 7347 -1130 7381
rect -1188 7332 -1130 7347
rect -930 7517 -872 7532
rect -930 7483 -918 7517
rect -884 7483 -872 7517
rect -930 7449 -872 7483
rect -930 7415 -918 7449
rect -884 7415 -872 7449
rect -930 7381 -872 7415
rect -930 7347 -918 7381
rect -884 7347 -872 7381
rect -930 7332 -872 7347
rect -672 7517 -614 7532
rect -672 7483 -660 7517
rect -626 7483 -614 7517
rect -672 7449 -614 7483
rect -672 7415 -660 7449
rect -626 7415 -614 7449
rect -672 7381 -614 7415
rect -672 7347 -660 7381
rect -626 7347 -614 7381
rect -672 7332 -614 7347
rect -414 7517 -356 7532
rect -414 7483 -402 7517
rect -368 7483 -356 7517
rect -414 7449 -356 7483
rect -414 7415 -402 7449
rect -368 7415 -356 7449
rect -414 7381 -356 7415
rect -414 7347 -402 7381
rect -368 7347 -356 7381
rect -414 7332 -356 7347
rect -156 7517 -98 7532
rect -156 7483 -144 7517
rect -110 7483 -98 7517
rect -156 7449 -98 7483
rect -156 7415 -144 7449
rect -110 7415 -98 7449
rect -156 7381 -98 7415
rect -156 7347 -144 7381
rect -110 7347 -98 7381
rect -156 7332 -98 7347
rect 102 7517 160 7532
rect 102 7483 114 7517
rect 148 7483 160 7517
rect 102 7449 160 7483
rect 102 7415 114 7449
rect 148 7415 160 7449
rect 102 7381 160 7415
rect 102 7347 114 7381
rect 148 7347 160 7381
rect 102 7332 160 7347
rect 360 7517 418 7532
rect 360 7483 372 7517
rect 406 7483 418 7517
rect 360 7449 418 7483
rect 360 7415 372 7449
rect 406 7415 418 7449
rect 360 7381 418 7415
rect 360 7347 372 7381
rect 406 7347 418 7381
rect 360 7332 418 7347
rect 618 7517 676 7532
rect 618 7483 630 7517
rect 664 7483 676 7517
rect 618 7449 676 7483
rect 618 7415 630 7449
rect 664 7415 676 7449
rect 618 7381 676 7415
rect 618 7347 630 7381
rect 664 7347 676 7381
rect 618 7332 676 7347
rect 876 7517 934 7532
rect 876 7483 888 7517
rect 922 7483 934 7517
rect 876 7449 934 7483
rect 876 7415 888 7449
rect 922 7415 934 7449
rect 876 7381 934 7415
rect 876 7347 888 7381
rect 922 7347 934 7381
rect 876 7332 934 7347
rect 1134 7517 1192 7532
rect 1134 7483 1146 7517
rect 1180 7483 1192 7517
rect 1134 7449 1192 7483
rect 1134 7415 1146 7449
rect 1180 7415 1192 7449
rect 1134 7381 1192 7415
rect 1134 7347 1146 7381
rect 1180 7347 1192 7381
rect 1134 7332 1192 7347
rect 1392 7517 1450 7532
rect 1392 7483 1404 7517
rect 1438 7483 1450 7517
rect 1392 7449 1450 7483
rect 1392 7415 1404 7449
rect 1438 7415 1450 7449
rect 1392 7381 1450 7415
rect 1392 7347 1404 7381
rect 1438 7347 1450 7381
rect 1392 7332 1450 7347
rect -2220 7099 -2162 7114
rect -2220 7065 -2208 7099
rect -2174 7065 -2162 7099
rect -2220 7031 -2162 7065
rect -2220 6997 -2208 7031
rect -2174 6997 -2162 7031
rect -2220 6963 -2162 6997
rect -2220 6929 -2208 6963
rect -2174 6929 -2162 6963
rect -2220 6914 -2162 6929
rect -1962 7099 -1904 7114
rect -1962 7065 -1950 7099
rect -1916 7065 -1904 7099
rect -1962 7031 -1904 7065
rect -1962 6997 -1950 7031
rect -1916 6997 -1904 7031
rect -1962 6963 -1904 6997
rect -1962 6929 -1950 6963
rect -1916 6929 -1904 6963
rect -1962 6914 -1904 6929
rect -1704 7099 -1646 7114
rect -1704 7065 -1692 7099
rect -1658 7065 -1646 7099
rect -1704 7031 -1646 7065
rect -1704 6997 -1692 7031
rect -1658 6997 -1646 7031
rect -1704 6963 -1646 6997
rect -1704 6929 -1692 6963
rect -1658 6929 -1646 6963
rect -1704 6914 -1646 6929
rect -1446 7099 -1388 7114
rect -1446 7065 -1434 7099
rect -1400 7065 -1388 7099
rect -1446 7031 -1388 7065
rect -1446 6997 -1434 7031
rect -1400 6997 -1388 7031
rect -1446 6963 -1388 6997
rect -1446 6929 -1434 6963
rect -1400 6929 -1388 6963
rect -1446 6914 -1388 6929
rect -1188 7099 -1130 7114
rect -1188 7065 -1176 7099
rect -1142 7065 -1130 7099
rect -1188 7031 -1130 7065
rect -1188 6997 -1176 7031
rect -1142 6997 -1130 7031
rect -1188 6963 -1130 6997
rect -1188 6929 -1176 6963
rect -1142 6929 -1130 6963
rect -1188 6914 -1130 6929
rect -930 7099 -872 7114
rect -930 7065 -918 7099
rect -884 7065 -872 7099
rect -930 7031 -872 7065
rect -930 6997 -918 7031
rect -884 6997 -872 7031
rect -930 6963 -872 6997
rect -930 6929 -918 6963
rect -884 6929 -872 6963
rect -930 6914 -872 6929
rect -672 7099 -614 7114
rect -672 7065 -660 7099
rect -626 7065 -614 7099
rect -672 7031 -614 7065
rect -672 6997 -660 7031
rect -626 6997 -614 7031
rect -672 6963 -614 6997
rect -672 6929 -660 6963
rect -626 6929 -614 6963
rect -672 6914 -614 6929
rect -414 7099 -356 7114
rect -414 7065 -402 7099
rect -368 7065 -356 7099
rect -414 7031 -356 7065
rect -414 6997 -402 7031
rect -368 6997 -356 7031
rect -414 6963 -356 6997
rect -414 6929 -402 6963
rect -368 6929 -356 6963
rect -414 6914 -356 6929
rect -156 7099 -98 7114
rect -156 7065 -144 7099
rect -110 7065 -98 7099
rect -156 7031 -98 7065
rect -156 6997 -144 7031
rect -110 6997 -98 7031
rect -156 6963 -98 6997
rect -156 6929 -144 6963
rect -110 6929 -98 6963
rect -156 6914 -98 6929
rect 102 7099 160 7114
rect 102 7065 114 7099
rect 148 7065 160 7099
rect 102 7031 160 7065
rect 102 6997 114 7031
rect 148 6997 160 7031
rect 102 6963 160 6997
rect 102 6929 114 6963
rect 148 6929 160 6963
rect 102 6914 160 6929
rect 360 7099 418 7114
rect 360 7065 372 7099
rect 406 7065 418 7099
rect 360 7031 418 7065
rect 360 6997 372 7031
rect 406 6997 418 7031
rect 360 6963 418 6997
rect 360 6929 372 6963
rect 406 6929 418 6963
rect 360 6914 418 6929
rect 618 7099 676 7114
rect 618 7065 630 7099
rect 664 7065 676 7099
rect 618 7031 676 7065
rect 618 6997 630 7031
rect 664 6997 676 7031
rect 618 6963 676 6997
rect 618 6929 630 6963
rect 664 6929 676 6963
rect 618 6914 676 6929
rect 876 7099 934 7114
rect 876 7065 888 7099
rect 922 7065 934 7099
rect 876 7031 934 7065
rect 876 6997 888 7031
rect 922 6997 934 7031
rect 876 6963 934 6997
rect 876 6929 888 6963
rect 922 6929 934 6963
rect 876 6914 934 6929
rect 1134 7099 1192 7114
rect 1134 7065 1146 7099
rect 1180 7065 1192 7099
rect 1134 7031 1192 7065
rect 1134 6997 1146 7031
rect 1180 6997 1192 7031
rect 1134 6963 1192 6997
rect 1134 6929 1146 6963
rect 1180 6929 1192 6963
rect 1134 6914 1192 6929
rect 1392 7099 1450 7114
rect 1392 7065 1404 7099
rect 1438 7065 1450 7099
rect 1392 7031 1450 7065
rect 1392 6997 1404 7031
rect 1438 6997 1450 7031
rect 1392 6963 1450 6997
rect 1392 6929 1404 6963
rect 1438 6929 1450 6963
rect 1392 6914 1450 6929
rect -2220 6681 -2162 6696
rect -2220 6647 -2208 6681
rect -2174 6647 -2162 6681
rect -2220 6613 -2162 6647
rect -2220 6579 -2208 6613
rect -2174 6579 -2162 6613
rect -2220 6545 -2162 6579
rect -2220 6511 -2208 6545
rect -2174 6511 -2162 6545
rect -2220 6496 -2162 6511
rect -1962 6681 -1904 6696
rect -1962 6647 -1950 6681
rect -1916 6647 -1904 6681
rect -1962 6613 -1904 6647
rect -1962 6579 -1950 6613
rect -1916 6579 -1904 6613
rect -1962 6545 -1904 6579
rect -1962 6511 -1950 6545
rect -1916 6511 -1904 6545
rect -1962 6496 -1904 6511
rect -1704 6681 -1646 6696
rect -1704 6647 -1692 6681
rect -1658 6647 -1646 6681
rect -1704 6613 -1646 6647
rect -1704 6579 -1692 6613
rect -1658 6579 -1646 6613
rect -1704 6545 -1646 6579
rect -1704 6511 -1692 6545
rect -1658 6511 -1646 6545
rect -1704 6496 -1646 6511
rect -1446 6681 -1388 6696
rect -1446 6647 -1434 6681
rect -1400 6647 -1388 6681
rect -1446 6613 -1388 6647
rect -1446 6579 -1434 6613
rect -1400 6579 -1388 6613
rect -1446 6545 -1388 6579
rect -1446 6511 -1434 6545
rect -1400 6511 -1388 6545
rect -1446 6496 -1388 6511
rect -1188 6681 -1130 6696
rect -1188 6647 -1176 6681
rect -1142 6647 -1130 6681
rect -1188 6613 -1130 6647
rect -1188 6579 -1176 6613
rect -1142 6579 -1130 6613
rect -1188 6545 -1130 6579
rect -1188 6511 -1176 6545
rect -1142 6511 -1130 6545
rect -1188 6496 -1130 6511
rect -930 6681 -872 6696
rect -930 6647 -918 6681
rect -884 6647 -872 6681
rect -930 6613 -872 6647
rect -930 6579 -918 6613
rect -884 6579 -872 6613
rect -930 6545 -872 6579
rect -930 6511 -918 6545
rect -884 6511 -872 6545
rect -930 6496 -872 6511
rect -672 6681 -614 6696
rect -672 6647 -660 6681
rect -626 6647 -614 6681
rect -672 6613 -614 6647
rect -672 6579 -660 6613
rect -626 6579 -614 6613
rect -672 6545 -614 6579
rect -672 6511 -660 6545
rect -626 6511 -614 6545
rect -672 6496 -614 6511
rect -414 6681 -356 6696
rect -414 6647 -402 6681
rect -368 6647 -356 6681
rect -414 6613 -356 6647
rect -414 6579 -402 6613
rect -368 6579 -356 6613
rect -414 6545 -356 6579
rect -414 6511 -402 6545
rect -368 6511 -356 6545
rect -414 6496 -356 6511
rect -156 6681 -98 6696
rect -156 6647 -144 6681
rect -110 6647 -98 6681
rect -156 6613 -98 6647
rect -156 6579 -144 6613
rect -110 6579 -98 6613
rect -156 6545 -98 6579
rect -156 6511 -144 6545
rect -110 6511 -98 6545
rect -156 6496 -98 6511
rect 102 6681 160 6696
rect 102 6647 114 6681
rect 148 6647 160 6681
rect 102 6613 160 6647
rect 102 6579 114 6613
rect 148 6579 160 6613
rect 102 6545 160 6579
rect 102 6511 114 6545
rect 148 6511 160 6545
rect 102 6496 160 6511
rect 360 6681 418 6696
rect 360 6647 372 6681
rect 406 6647 418 6681
rect 360 6613 418 6647
rect 360 6579 372 6613
rect 406 6579 418 6613
rect 360 6545 418 6579
rect 360 6511 372 6545
rect 406 6511 418 6545
rect 360 6496 418 6511
rect 618 6681 676 6696
rect 618 6647 630 6681
rect 664 6647 676 6681
rect 618 6613 676 6647
rect 618 6579 630 6613
rect 664 6579 676 6613
rect 618 6545 676 6579
rect 618 6511 630 6545
rect 664 6511 676 6545
rect 618 6496 676 6511
rect 876 6681 934 6696
rect 876 6647 888 6681
rect 922 6647 934 6681
rect 876 6613 934 6647
rect 876 6579 888 6613
rect 922 6579 934 6613
rect 876 6545 934 6579
rect 876 6511 888 6545
rect 922 6511 934 6545
rect 876 6496 934 6511
rect 1134 6681 1192 6696
rect 1134 6647 1146 6681
rect 1180 6647 1192 6681
rect 1134 6613 1192 6647
rect 1134 6579 1146 6613
rect 1180 6579 1192 6613
rect 1134 6545 1192 6579
rect 1134 6511 1146 6545
rect 1180 6511 1192 6545
rect 1134 6496 1192 6511
rect 1392 6681 1450 6696
rect 1392 6647 1404 6681
rect 1438 6647 1450 6681
rect 1392 6613 1450 6647
rect 1392 6579 1404 6613
rect 1438 6579 1450 6613
rect 1392 6545 1450 6579
rect 1392 6511 1404 6545
rect 1438 6511 1450 6545
rect 1392 6496 1450 6511
rect -2220 6263 -2162 6278
rect -2220 6229 -2208 6263
rect -2174 6229 -2162 6263
rect -2220 6195 -2162 6229
rect -2220 6161 -2208 6195
rect -2174 6161 -2162 6195
rect -2220 6127 -2162 6161
rect -2220 6093 -2208 6127
rect -2174 6093 -2162 6127
rect -2220 6078 -2162 6093
rect -1962 6263 -1904 6278
rect -1962 6229 -1950 6263
rect -1916 6229 -1904 6263
rect -1962 6195 -1904 6229
rect -1962 6161 -1950 6195
rect -1916 6161 -1904 6195
rect -1962 6127 -1904 6161
rect -1962 6093 -1950 6127
rect -1916 6093 -1904 6127
rect -1962 6078 -1904 6093
rect -1704 6263 -1646 6278
rect -1704 6229 -1692 6263
rect -1658 6229 -1646 6263
rect -1704 6195 -1646 6229
rect -1704 6161 -1692 6195
rect -1658 6161 -1646 6195
rect -1704 6127 -1646 6161
rect -1704 6093 -1692 6127
rect -1658 6093 -1646 6127
rect -1704 6078 -1646 6093
rect -1446 6263 -1388 6278
rect -1446 6229 -1434 6263
rect -1400 6229 -1388 6263
rect -1446 6195 -1388 6229
rect -1446 6161 -1434 6195
rect -1400 6161 -1388 6195
rect -1446 6127 -1388 6161
rect -1446 6093 -1434 6127
rect -1400 6093 -1388 6127
rect -1446 6078 -1388 6093
rect -1188 6263 -1130 6278
rect -1188 6229 -1176 6263
rect -1142 6229 -1130 6263
rect -1188 6195 -1130 6229
rect -1188 6161 -1176 6195
rect -1142 6161 -1130 6195
rect -1188 6127 -1130 6161
rect -1188 6093 -1176 6127
rect -1142 6093 -1130 6127
rect -1188 6078 -1130 6093
rect -930 6263 -872 6278
rect -930 6229 -918 6263
rect -884 6229 -872 6263
rect -930 6195 -872 6229
rect -930 6161 -918 6195
rect -884 6161 -872 6195
rect -930 6127 -872 6161
rect -930 6093 -918 6127
rect -884 6093 -872 6127
rect -930 6078 -872 6093
rect -672 6263 -614 6278
rect -672 6229 -660 6263
rect -626 6229 -614 6263
rect -672 6195 -614 6229
rect -672 6161 -660 6195
rect -626 6161 -614 6195
rect -672 6127 -614 6161
rect -672 6093 -660 6127
rect -626 6093 -614 6127
rect -672 6078 -614 6093
rect -414 6263 -356 6278
rect -414 6229 -402 6263
rect -368 6229 -356 6263
rect -414 6195 -356 6229
rect -414 6161 -402 6195
rect -368 6161 -356 6195
rect -414 6127 -356 6161
rect -414 6093 -402 6127
rect -368 6093 -356 6127
rect -414 6078 -356 6093
rect -156 6263 -98 6278
rect -156 6229 -144 6263
rect -110 6229 -98 6263
rect -156 6195 -98 6229
rect -156 6161 -144 6195
rect -110 6161 -98 6195
rect -156 6127 -98 6161
rect -156 6093 -144 6127
rect -110 6093 -98 6127
rect -156 6078 -98 6093
rect 102 6263 160 6278
rect 102 6229 114 6263
rect 148 6229 160 6263
rect 102 6195 160 6229
rect 102 6161 114 6195
rect 148 6161 160 6195
rect 102 6127 160 6161
rect 102 6093 114 6127
rect 148 6093 160 6127
rect 102 6078 160 6093
rect 360 6263 418 6278
rect 360 6229 372 6263
rect 406 6229 418 6263
rect 360 6195 418 6229
rect 360 6161 372 6195
rect 406 6161 418 6195
rect 360 6127 418 6161
rect 360 6093 372 6127
rect 406 6093 418 6127
rect 360 6078 418 6093
rect 618 6263 676 6278
rect 618 6229 630 6263
rect 664 6229 676 6263
rect 618 6195 676 6229
rect 618 6161 630 6195
rect 664 6161 676 6195
rect 618 6127 676 6161
rect 618 6093 630 6127
rect 664 6093 676 6127
rect 618 6078 676 6093
rect 876 6263 934 6278
rect 876 6229 888 6263
rect 922 6229 934 6263
rect 876 6195 934 6229
rect 876 6161 888 6195
rect 922 6161 934 6195
rect 876 6127 934 6161
rect 876 6093 888 6127
rect 922 6093 934 6127
rect 876 6078 934 6093
rect 1134 6263 1192 6278
rect 1134 6229 1146 6263
rect 1180 6229 1192 6263
rect 1134 6195 1192 6229
rect 1134 6161 1146 6195
rect 1180 6161 1192 6195
rect 1134 6127 1192 6161
rect 1134 6093 1146 6127
rect 1180 6093 1192 6127
rect 1134 6078 1192 6093
rect 1392 6263 1450 6278
rect 1392 6229 1404 6263
rect 1438 6229 1450 6263
rect 1392 6195 1450 6229
rect 1392 6161 1404 6195
rect 1438 6161 1450 6195
rect 1392 6127 1450 6161
rect 1392 6093 1404 6127
rect 1438 6093 1450 6127
rect 1392 6078 1450 6093
rect -2220 5845 -2162 5860
rect -2220 5811 -2208 5845
rect -2174 5811 -2162 5845
rect -2220 5777 -2162 5811
rect -2220 5743 -2208 5777
rect -2174 5743 -2162 5777
rect -2220 5709 -2162 5743
rect -2220 5675 -2208 5709
rect -2174 5675 -2162 5709
rect -2220 5660 -2162 5675
rect -1962 5845 -1904 5860
rect -1962 5811 -1950 5845
rect -1916 5811 -1904 5845
rect -1962 5777 -1904 5811
rect -1962 5743 -1950 5777
rect -1916 5743 -1904 5777
rect -1962 5709 -1904 5743
rect -1962 5675 -1950 5709
rect -1916 5675 -1904 5709
rect -1962 5660 -1904 5675
rect -1704 5845 -1646 5860
rect -1704 5811 -1692 5845
rect -1658 5811 -1646 5845
rect -1704 5777 -1646 5811
rect -1704 5743 -1692 5777
rect -1658 5743 -1646 5777
rect -1704 5709 -1646 5743
rect -1704 5675 -1692 5709
rect -1658 5675 -1646 5709
rect -1704 5660 -1646 5675
rect -1446 5845 -1388 5860
rect -1446 5811 -1434 5845
rect -1400 5811 -1388 5845
rect -1446 5777 -1388 5811
rect -1446 5743 -1434 5777
rect -1400 5743 -1388 5777
rect -1446 5709 -1388 5743
rect -1446 5675 -1434 5709
rect -1400 5675 -1388 5709
rect -1446 5660 -1388 5675
rect -1188 5845 -1130 5860
rect -1188 5811 -1176 5845
rect -1142 5811 -1130 5845
rect -1188 5777 -1130 5811
rect -1188 5743 -1176 5777
rect -1142 5743 -1130 5777
rect -1188 5709 -1130 5743
rect -1188 5675 -1176 5709
rect -1142 5675 -1130 5709
rect -1188 5660 -1130 5675
rect -930 5845 -872 5860
rect -930 5811 -918 5845
rect -884 5811 -872 5845
rect -930 5777 -872 5811
rect -930 5743 -918 5777
rect -884 5743 -872 5777
rect -930 5709 -872 5743
rect -930 5675 -918 5709
rect -884 5675 -872 5709
rect -930 5660 -872 5675
rect -672 5845 -614 5860
rect -672 5811 -660 5845
rect -626 5811 -614 5845
rect -672 5777 -614 5811
rect -672 5743 -660 5777
rect -626 5743 -614 5777
rect -672 5709 -614 5743
rect -672 5675 -660 5709
rect -626 5675 -614 5709
rect -672 5660 -614 5675
rect -414 5845 -356 5860
rect -414 5811 -402 5845
rect -368 5811 -356 5845
rect -414 5777 -356 5811
rect -414 5743 -402 5777
rect -368 5743 -356 5777
rect -414 5709 -356 5743
rect -414 5675 -402 5709
rect -368 5675 -356 5709
rect -414 5660 -356 5675
rect -156 5845 -98 5860
rect -156 5811 -144 5845
rect -110 5811 -98 5845
rect -156 5777 -98 5811
rect -156 5743 -144 5777
rect -110 5743 -98 5777
rect -156 5709 -98 5743
rect -156 5675 -144 5709
rect -110 5675 -98 5709
rect -156 5660 -98 5675
rect 102 5845 160 5860
rect 102 5811 114 5845
rect 148 5811 160 5845
rect 102 5777 160 5811
rect 102 5743 114 5777
rect 148 5743 160 5777
rect 102 5709 160 5743
rect 102 5675 114 5709
rect 148 5675 160 5709
rect 102 5660 160 5675
rect 360 5845 418 5860
rect 360 5811 372 5845
rect 406 5811 418 5845
rect 360 5777 418 5811
rect 360 5743 372 5777
rect 406 5743 418 5777
rect 360 5709 418 5743
rect 360 5675 372 5709
rect 406 5675 418 5709
rect 360 5660 418 5675
rect 618 5845 676 5860
rect 618 5811 630 5845
rect 664 5811 676 5845
rect 618 5777 676 5811
rect 618 5743 630 5777
rect 664 5743 676 5777
rect 618 5709 676 5743
rect 618 5675 630 5709
rect 664 5675 676 5709
rect 618 5660 676 5675
rect 876 5845 934 5860
rect 876 5811 888 5845
rect 922 5811 934 5845
rect 876 5777 934 5811
rect 876 5743 888 5777
rect 922 5743 934 5777
rect 876 5709 934 5743
rect 876 5675 888 5709
rect 922 5675 934 5709
rect 876 5660 934 5675
rect 1134 5845 1192 5860
rect 1134 5811 1146 5845
rect 1180 5811 1192 5845
rect 1134 5777 1192 5811
rect 1134 5743 1146 5777
rect 1180 5743 1192 5777
rect 1134 5709 1192 5743
rect 1134 5675 1146 5709
rect 1180 5675 1192 5709
rect 1134 5660 1192 5675
rect 1392 5845 1450 5860
rect 1392 5811 1404 5845
rect 1438 5811 1450 5845
rect 1392 5777 1450 5811
rect 1392 5743 1404 5777
rect 1438 5743 1450 5777
rect 1392 5709 1450 5743
rect 1392 5675 1404 5709
rect 1438 5675 1450 5709
rect 1392 5660 1450 5675
rect -2220 5427 -2162 5442
rect -2220 5393 -2208 5427
rect -2174 5393 -2162 5427
rect -2220 5359 -2162 5393
rect -2220 5325 -2208 5359
rect -2174 5325 -2162 5359
rect -2220 5291 -2162 5325
rect -2220 5257 -2208 5291
rect -2174 5257 -2162 5291
rect -2220 5242 -2162 5257
rect -1962 5427 -1904 5442
rect -1962 5393 -1950 5427
rect -1916 5393 -1904 5427
rect -1962 5359 -1904 5393
rect -1962 5325 -1950 5359
rect -1916 5325 -1904 5359
rect -1962 5291 -1904 5325
rect -1962 5257 -1950 5291
rect -1916 5257 -1904 5291
rect -1962 5242 -1904 5257
rect -1704 5427 -1646 5442
rect -1704 5393 -1692 5427
rect -1658 5393 -1646 5427
rect -1704 5359 -1646 5393
rect -1704 5325 -1692 5359
rect -1658 5325 -1646 5359
rect -1704 5291 -1646 5325
rect -1704 5257 -1692 5291
rect -1658 5257 -1646 5291
rect -1704 5242 -1646 5257
rect -1446 5427 -1388 5442
rect -1446 5393 -1434 5427
rect -1400 5393 -1388 5427
rect -1446 5359 -1388 5393
rect -1446 5325 -1434 5359
rect -1400 5325 -1388 5359
rect -1446 5291 -1388 5325
rect -1446 5257 -1434 5291
rect -1400 5257 -1388 5291
rect -1446 5242 -1388 5257
rect -1188 5427 -1130 5442
rect -1188 5393 -1176 5427
rect -1142 5393 -1130 5427
rect -1188 5359 -1130 5393
rect -1188 5325 -1176 5359
rect -1142 5325 -1130 5359
rect -1188 5291 -1130 5325
rect -1188 5257 -1176 5291
rect -1142 5257 -1130 5291
rect -1188 5242 -1130 5257
rect -930 5427 -872 5442
rect -930 5393 -918 5427
rect -884 5393 -872 5427
rect -930 5359 -872 5393
rect -930 5325 -918 5359
rect -884 5325 -872 5359
rect -930 5291 -872 5325
rect -930 5257 -918 5291
rect -884 5257 -872 5291
rect -930 5242 -872 5257
rect -672 5427 -614 5442
rect -672 5393 -660 5427
rect -626 5393 -614 5427
rect -672 5359 -614 5393
rect -672 5325 -660 5359
rect -626 5325 -614 5359
rect -672 5291 -614 5325
rect -672 5257 -660 5291
rect -626 5257 -614 5291
rect -672 5242 -614 5257
rect -414 5427 -356 5442
rect -414 5393 -402 5427
rect -368 5393 -356 5427
rect -414 5359 -356 5393
rect -414 5325 -402 5359
rect -368 5325 -356 5359
rect -414 5291 -356 5325
rect -414 5257 -402 5291
rect -368 5257 -356 5291
rect -414 5242 -356 5257
rect -156 5427 -98 5442
rect -156 5393 -144 5427
rect -110 5393 -98 5427
rect -156 5359 -98 5393
rect -156 5325 -144 5359
rect -110 5325 -98 5359
rect -156 5291 -98 5325
rect -156 5257 -144 5291
rect -110 5257 -98 5291
rect -156 5242 -98 5257
rect 102 5427 160 5442
rect 102 5393 114 5427
rect 148 5393 160 5427
rect 102 5359 160 5393
rect 102 5325 114 5359
rect 148 5325 160 5359
rect 102 5291 160 5325
rect 102 5257 114 5291
rect 148 5257 160 5291
rect 102 5242 160 5257
rect 360 5427 418 5442
rect 360 5393 372 5427
rect 406 5393 418 5427
rect 360 5359 418 5393
rect 360 5325 372 5359
rect 406 5325 418 5359
rect 360 5291 418 5325
rect 360 5257 372 5291
rect 406 5257 418 5291
rect 360 5242 418 5257
rect 618 5427 676 5442
rect 618 5393 630 5427
rect 664 5393 676 5427
rect 618 5359 676 5393
rect 618 5325 630 5359
rect 664 5325 676 5359
rect 618 5291 676 5325
rect 618 5257 630 5291
rect 664 5257 676 5291
rect 618 5242 676 5257
rect 876 5427 934 5442
rect 876 5393 888 5427
rect 922 5393 934 5427
rect 876 5359 934 5393
rect 876 5325 888 5359
rect 922 5325 934 5359
rect 876 5291 934 5325
rect 876 5257 888 5291
rect 922 5257 934 5291
rect 876 5242 934 5257
rect 1134 5427 1192 5442
rect 1134 5393 1146 5427
rect 1180 5393 1192 5427
rect 1134 5359 1192 5393
rect 1134 5325 1146 5359
rect 1180 5325 1192 5359
rect 1134 5291 1192 5325
rect 1134 5257 1146 5291
rect 1180 5257 1192 5291
rect 1134 5242 1192 5257
rect 1392 5427 1450 5442
rect 1392 5393 1404 5427
rect 1438 5393 1450 5427
rect 1392 5359 1450 5393
rect 1392 5325 1404 5359
rect 1438 5325 1450 5359
rect 1392 5291 1450 5325
rect 1392 5257 1404 5291
rect 1438 5257 1450 5291
rect 1392 5242 1450 5257
rect -2220 5009 -2162 5024
rect -2220 4975 -2208 5009
rect -2174 4975 -2162 5009
rect -2220 4941 -2162 4975
rect -2220 4907 -2208 4941
rect -2174 4907 -2162 4941
rect -2220 4873 -2162 4907
rect -2220 4839 -2208 4873
rect -2174 4839 -2162 4873
rect -2220 4824 -2162 4839
rect -1962 5009 -1904 5024
rect -1962 4975 -1950 5009
rect -1916 4975 -1904 5009
rect -1962 4941 -1904 4975
rect -1962 4907 -1950 4941
rect -1916 4907 -1904 4941
rect -1962 4873 -1904 4907
rect -1962 4839 -1950 4873
rect -1916 4839 -1904 4873
rect -1962 4824 -1904 4839
rect -1704 5009 -1646 5024
rect -1704 4975 -1692 5009
rect -1658 4975 -1646 5009
rect -1704 4941 -1646 4975
rect -1704 4907 -1692 4941
rect -1658 4907 -1646 4941
rect -1704 4873 -1646 4907
rect -1704 4839 -1692 4873
rect -1658 4839 -1646 4873
rect -1704 4824 -1646 4839
rect -1446 5009 -1388 5024
rect -1446 4975 -1434 5009
rect -1400 4975 -1388 5009
rect -1446 4941 -1388 4975
rect -1446 4907 -1434 4941
rect -1400 4907 -1388 4941
rect -1446 4873 -1388 4907
rect -1446 4839 -1434 4873
rect -1400 4839 -1388 4873
rect -1446 4824 -1388 4839
rect -1188 5009 -1130 5024
rect -1188 4975 -1176 5009
rect -1142 4975 -1130 5009
rect -1188 4941 -1130 4975
rect -1188 4907 -1176 4941
rect -1142 4907 -1130 4941
rect -1188 4873 -1130 4907
rect -1188 4839 -1176 4873
rect -1142 4839 -1130 4873
rect -1188 4824 -1130 4839
rect -930 5009 -872 5024
rect -930 4975 -918 5009
rect -884 4975 -872 5009
rect -930 4941 -872 4975
rect -930 4907 -918 4941
rect -884 4907 -872 4941
rect -930 4873 -872 4907
rect -930 4839 -918 4873
rect -884 4839 -872 4873
rect -930 4824 -872 4839
rect -672 5009 -614 5024
rect -672 4975 -660 5009
rect -626 4975 -614 5009
rect -672 4941 -614 4975
rect -672 4907 -660 4941
rect -626 4907 -614 4941
rect -672 4873 -614 4907
rect -672 4839 -660 4873
rect -626 4839 -614 4873
rect -672 4824 -614 4839
rect -414 5009 -356 5024
rect -414 4975 -402 5009
rect -368 4975 -356 5009
rect -414 4941 -356 4975
rect -414 4907 -402 4941
rect -368 4907 -356 4941
rect -414 4873 -356 4907
rect -414 4839 -402 4873
rect -368 4839 -356 4873
rect -414 4824 -356 4839
rect -156 5009 -98 5024
rect -156 4975 -144 5009
rect -110 4975 -98 5009
rect -156 4941 -98 4975
rect -156 4907 -144 4941
rect -110 4907 -98 4941
rect -156 4873 -98 4907
rect -156 4839 -144 4873
rect -110 4839 -98 4873
rect -156 4824 -98 4839
rect 102 5009 160 5024
rect 102 4975 114 5009
rect 148 4975 160 5009
rect 102 4941 160 4975
rect 102 4907 114 4941
rect 148 4907 160 4941
rect 102 4873 160 4907
rect 102 4839 114 4873
rect 148 4839 160 4873
rect 102 4824 160 4839
rect 360 5009 418 5024
rect 360 4975 372 5009
rect 406 4975 418 5009
rect 360 4941 418 4975
rect 360 4907 372 4941
rect 406 4907 418 4941
rect 360 4873 418 4907
rect 360 4839 372 4873
rect 406 4839 418 4873
rect 360 4824 418 4839
rect 618 5009 676 5024
rect 618 4975 630 5009
rect 664 4975 676 5009
rect 618 4941 676 4975
rect 618 4907 630 4941
rect 664 4907 676 4941
rect 618 4873 676 4907
rect 618 4839 630 4873
rect 664 4839 676 4873
rect 618 4824 676 4839
rect 876 5009 934 5024
rect 876 4975 888 5009
rect 922 4975 934 5009
rect 876 4941 934 4975
rect 876 4907 888 4941
rect 922 4907 934 4941
rect 876 4873 934 4907
rect 876 4839 888 4873
rect 922 4839 934 4873
rect 876 4824 934 4839
rect 1134 5009 1192 5024
rect 1134 4975 1146 5009
rect 1180 4975 1192 5009
rect 1134 4941 1192 4975
rect 1134 4907 1146 4941
rect 1180 4907 1192 4941
rect 1134 4873 1192 4907
rect 1134 4839 1146 4873
rect 1180 4839 1192 4873
rect 1134 4824 1192 4839
rect 1392 5009 1450 5024
rect 1392 4975 1404 5009
rect 1438 4975 1450 5009
rect 1392 4941 1450 4975
rect 1392 4907 1404 4941
rect 1438 4907 1450 4941
rect 1392 4873 1450 4907
rect 1392 4839 1404 4873
rect 1438 4839 1450 4873
rect 1392 4824 1450 4839
rect -2220 4591 -2162 4606
rect -2220 4557 -2208 4591
rect -2174 4557 -2162 4591
rect -2220 4523 -2162 4557
rect -2220 4489 -2208 4523
rect -2174 4489 -2162 4523
rect -2220 4455 -2162 4489
rect -2220 4421 -2208 4455
rect -2174 4421 -2162 4455
rect -2220 4406 -2162 4421
rect -1962 4591 -1904 4606
rect -1962 4557 -1950 4591
rect -1916 4557 -1904 4591
rect -1962 4523 -1904 4557
rect -1962 4489 -1950 4523
rect -1916 4489 -1904 4523
rect -1962 4455 -1904 4489
rect -1962 4421 -1950 4455
rect -1916 4421 -1904 4455
rect -1962 4406 -1904 4421
rect -1704 4591 -1646 4606
rect -1704 4557 -1692 4591
rect -1658 4557 -1646 4591
rect -1704 4523 -1646 4557
rect -1704 4489 -1692 4523
rect -1658 4489 -1646 4523
rect -1704 4455 -1646 4489
rect -1704 4421 -1692 4455
rect -1658 4421 -1646 4455
rect -1704 4406 -1646 4421
rect -1446 4591 -1388 4606
rect -1446 4557 -1434 4591
rect -1400 4557 -1388 4591
rect -1446 4523 -1388 4557
rect -1446 4489 -1434 4523
rect -1400 4489 -1388 4523
rect -1446 4455 -1388 4489
rect -1446 4421 -1434 4455
rect -1400 4421 -1388 4455
rect -1446 4406 -1388 4421
rect -1188 4591 -1130 4606
rect -1188 4557 -1176 4591
rect -1142 4557 -1130 4591
rect -1188 4523 -1130 4557
rect -1188 4489 -1176 4523
rect -1142 4489 -1130 4523
rect -1188 4455 -1130 4489
rect -1188 4421 -1176 4455
rect -1142 4421 -1130 4455
rect -1188 4406 -1130 4421
rect -930 4591 -872 4606
rect -930 4557 -918 4591
rect -884 4557 -872 4591
rect -930 4523 -872 4557
rect -930 4489 -918 4523
rect -884 4489 -872 4523
rect -930 4455 -872 4489
rect -930 4421 -918 4455
rect -884 4421 -872 4455
rect -930 4406 -872 4421
rect -672 4591 -614 4606
rect -672 4557 -660 4591
rect -626 4557 -614 4591
rect -672 4523 -614 4557
rect -672 4489 -660 4523
rect -626 4489 -614 4523
rect -672 4455 -614 4489
rect -672 4421 -660 4455
rect -626 4421 -614 4455
rect -672 4406 -614 4421
rect -414 4591 -356 4606
rect -414 4557 -402 4591
rect -368 4557 -356 4591
rect -414 4523 -356 4557
rect -414 4489 -402 4523
rect -368 4489 -356 4523
rect -414 4455 -356 4489
rect -414 4421 -402 4455
rect -368 4421 -356 4455
rect -414 4406 -356 4421
rect -156 4591 -98 4606
rect -156 4557 -144 4591
rect -110 4557 -98 4591
rect -156 4523 -98 4557
rect -156 4489 -144 4523
rect -110 4489 -98 4523
rect -156 4455 -98 4489
rect -156 4421 -144 4455
rect -110 4421 -98 4455
rect -156 4406 -98 4421
rect 102 4591 160 4606
rect 102 4557 114 4591
rect 148 4557 160 4591
rect 102 4523 160 4557
rect 102 4489 114 4523
rect 148 4489 160 4523
rect 102 4455 160 4489
rect 102 4421 114 4455
rect 148 4421 160 4455
rect 102 4406 160 4421
rect 360 4591 418 4606
rect 360 4557 372 4591
rect 406 4557 418 4591
rect 360 4523 418 4557
rect 360 4489 372 4523
rect 406 4489 418 4523
rect 360 4455 418 4489
rect 360 4421 372 4455
rect 406 4421 418 4455
rect 360 4406 418 4421
rect 618 4591 676 4606
rect 618 4557 630 4591
rect 664 4557 676 4591
rect 618 4523 676 4557
rect 618 4489 630 4523
rect 664 4489 676 4523
rect 618 4455 676 4489
rect 618 4421 630 4455
rect 664 4421 676 4455
rect 618 4406 676 4421
rect 876 4591 934 4606
rect 876 4557 888 4591
rect 922 4557 934 4591
rect 876 4523 934 4557
rect 876 4489 888 4523
rect 922 4489 934 4523
rect 876 4455 934 4489
rect 876 4421 888 4455
rect 922 4421 934 4455
rect 876 4406 934 4421
rect 1134 4591 1192 4606
rect 1134 4557 1146 4591
rect 1180 4557 1192 4591
rect 1134 4523 1192 4557
rect 1134 4489 1146 4523
rect 1180 4489 1192 4523
rect 1134 4455 1192 4489
rect 1134 4421 1146 4455
rect 1180 4421 1192 4455
rect 1134 4406 1192 4421
rect 1392 4591 1450 4606
rect 1392 4557 1404 4591
rect 1438 4557 1450 4591
rect 1392 4523 1450 4557
rect 1392 4489 1404 4523
rect 1438 4489 1450 4523
rect 1392 4455 1450 4489
rect 1392 4421 1404 4455
rect 1438 4421 1450 4455
rect 1392 4406 1450 4421
rect -2220 4173 -2162 4188
rect -2220 4139 -2208 4173
rect -2174 4139 -2162 4173
rect -2220 4105 -2162 4139
rect -2220 4071 -2208 4105
rect -2174 4071 -2162 4105
rect -2220 4037 -2162 4071
rect -2220 4003 -2208 4037
rect -2174 4003 -2162 4037
rect -2220 3988 -2162 4003
rect -1962 4173 -1904 4188
rect -1962 4139 -1950 4173
rect -1916 4139 -1904 4173
rect -1962 4105 -1904 4139
rect -1962 4071 -1950 4105
rect -1916 4071 -1904 4105
rect -1962 4037 -1904 4071
rect -1962 4003 -1950 4037
rect -1916 4003 -1904 4037
rect -1962 3988 -1904 4003
rect -1704 4173 -1646 4188
rect -1704 4139 -1692 4173
rect -1658 4139 -1646 4173
rect -1704 4105 -1646 4139
rect -1704 4071 -1692 4105
rect -1658 4071 -1646 4105
rect -1704 4037 -1646 4071
rect -1704 4003 -1692 4037
rect -1658 4003 -1646 4037
rect -1704 3988 -1646 4003
rect -1446 4173 -1388 4188
rect -1446 4139 -1434 4173
rect -1400 4139 -1388 4173
rect -1446 4105 -1388 4139
rect -1446 4071 -1434 4105
rect -1400 4071 -1388 4105
rect -1446 4037 -1388 4071
rect -1446 4003 -1434 4037
rect -1400 4003 -1388 4037
rect -1446 3988 -1388 4003
rect -1188 4173 -1130 4188
rect -1188 4139 -1176 4173
rect -1142 4139 -1130 4173
rect -1188 4105 -1130 4139
rect -1188 4071 -1176 4105
rect -1142 4071 -1130 4105
rect -1188 4037 -1130 4071
rect -1188 4003 -1176 4037
rect -1142 4003 -1130 4037
rect -1188 3988 -1130 4003
rect -930 4173 -872 4188
rect -930 4139 -918 4173
rect -884 4139 -872 4173
rect -930 4105 -872 4139
rect -930 4071 -918 4105
rect -884 4071 -872 4105
rect -930 4037 -872 4071
rect -930 4003 -918 4037
rect -884 4003 -872 4037
rect -930 3988 -872 4003
rect -672 4173 -614 4188
rect -672 4139 -660 4173
rect -626 4139 -614 4173
rect -672 4105 -614 4139
rect -672 4071 -660 4105
rect -626 4071 -614 4105
rect -672 4037 -614 4071
rect -672 4003 -660 4037
rect -626 4003 -614 4037
rect -672 3988 -614 4003
rect -414 4173 -356 4188
rect -414 4139 -402 4173
rect -368 4139 -356 4173
rect -414 4105 -356 4139
rect -414 4071 -402 4105
rect -368 4071 -356 4105
rect -414 4037 -356 4071
rect -414 4003 -402 4037
rect -368 4003 -356 4037
rect -414 3988 -356 4003
rect -156 4173 -98 4188
rect -156 4139 -144 4173
rect -110 4139 -98 4173
rect -156 4105 -98 4139
rect -156 4071 -144 4105
rect -110 4071 -98 4105
rect -156 4037 -98 4071
rect -156 4003 -144 4037
rect -110 4003 -98 4037
rect -156 3988 -98 4003
rect 102 4173 160 4188
rect 102 4139 114 4173
rect 148 4139 160 4173
rect 102 4105 160 4139
rect 102 4071 114 4105
rect 148 4071 160 4105
rect 102 4037 160 4071
rect 102 4003 114 4037
rect 148 4003 160 4037
rect 102 3988 160 4003
rect 360 4173 418 4188
rect 360 4139 372 4173
rect 406 4139 418 4173
rect 360 4105 418 4139
rect 360 4071 372 4105
rect 406 4071 418 4105
rect 360 4037 418 4071
rect 360 4003 372 4037
rect 406 4003 418 4037
rect 360 3988 418 4003
rect 618 4173 676 4188
rect 618 4139 630 4173
rect 664 4139 676 4173
rect 618 4105 676 4139
rect 618 4071 630 4105
rect 664 4071 676 4105
rect 618 4037 676 4071
rect 618 4003 630 4037
rect 664 4003 676 4037
rect 618 3988 676 4003
rect 876 4173 934 4188
rect 876 4139 888 4173
rect 922 4139 934 4173
rect 876 4105 934 4139
rect 876 4071 888 4105
rect 922 4071 934 4105
rect 876 4037 934 4071
rect 876 4003 888 4037
rect 922 4003 934 4037
rect 876 3988 934 4003
rect 1134 4173 1192 4188
rect 1134 4139 1146 4173
rect 1180 4139 1192 4173
rect 1134 4105 1192 4139
rect 1134 4071 1146 4105
rect 1180 4071 1192 4105
rect 1134 4037 1192 4071
rect 1134 4003 1146 4037
rect 1180 4003 1192 4037
rect 1134 3988 1192 4003
rect 1392 4173 1450 4188
rect 1392 4139 1404 4173
rect 1438 4139 1450 4173
rect 1392 4105 1450 4139
rect 1392 4071 1404 4105
rect 1438 4071 1450 4105
rect 1392 4037 1450 4071
rect 1392 4003 1404 4037
rect 1438 4003 1450 4037
rect 1392 3988 1450 4003
rect 3610 7296 3668 7311
rect 3610 7262 3622 7296
rect 3656 7262 3668 7296
rect 3610 7228 3668 7262
rect 3610 7194 3622 7228
rect 3656 7194 3668 7228
rect 3610 7160 3668 7194
rect 3610 7126 3622 7160
rect 3656 7126 3668 7160
rect 3610 7111 3668 7126
rect 3868 7296 3926 7311
rect 3868 7262 3880 7296
rect 3914 7262 3926 7296
rect 3868 7228 3926 7262
rect 3868 7194 3880 7228
rect 3914 7194 3926 7228
rect 3868 7160 3926 7194
rect 3868 7126 3880 7160
rect 3914 7126 3926 7160
rect 3868 7111 3926 7126
rect 4126 7296 4184 7311
rect 4126 7262 4138 7296
rect 4172 7262 4184 7296
rect 4126 7228 4184 7262
rect 4126 7194 4138 7228
rect 4172 7194 4184 7228
rect 4126 7160 4184 7194
rect 4126 7126 4138 7160
rect 4172 7126 4184 7160
rect 4126 7111 4184 7126
rect 4384 7296 4442 7311
rect 4384 7262 4396 7296
rect 4430 7262 4442 7296
rect 4384 7228 4442 7262
rect 4384 7194 4396 7228
rect 4430 7194 4442 7228
rect 4384 7160 4442 7194
rect 4384 7126 4396 7160
rect 4430 7126 4442 7160
rect 4384 7111 4442 7126
rect 4642 7296 4700 7311
rect 4642 7262 4654 7296
rect 4688 7262 4700 7296
rect 4642 7228 4700 7262
rect 4642 7194 4654 7228
rect 4688 7194 4700 7228
rect 4642 7160 4700 7194
rect 4642 7126 4654 7160
rect 4688 7126 4700 7160
rect 4642 7111 4700 7126
rect 4900 7296 4958 7311
rect 4900 7262 4912 7296
rect 4946 7262 4958 7296
rect 4900 7228 4958 7262
rect 4900 7194 4912 7228
rect 4946 7194 4958 7228
rect 4900 7160 4958 7194
rect 4900 7126 4912 7160
rect 4946 7126 4958 7160
rect 4900 7111 4958 7126
rect 5158 7296 5216 7311
rect 5158 7262 5170 7296
rect 5204 7262 5216 7296
rect 5158 7228 5216 7262
rect 5158 7194 5170 7228
rect 5204 7194 5216 7228
rect 5158 7160 5216 7194
rect 5158 7126 5170 7160
rect 5204 7126 5216 7160
rect 5158 7111 5216 7126
rect 5416 7296 5474 7311
rect 5416 7262 5428 7296
rect 5462 7262 5474 7296
rect 5416 7228 5474 7262
rect 5416 7194 5428 7228
rect 5462 7194 5474 7228
rect 5416 7160 5474 7194
rect 5416 7126 5428 7160
rect 5462 7126 5474 7160
rect 5416 7111 5474 7126
rect 5674 7296 5732 7311
rect 5674 7262 5686 7296
rect 5720 7262 5732 7296
rect 5674 7228 5732 7262
rect 5674 7194 5686 7228
rect 5720 7194 5732 7228
rect 5674 7160 5732 7194
rect 5674 7126 5686 7160
rect 5720 7126 5732 7160
rect 5674 7111 5732 7126
rect 5932 7296 5990 7311
rect 5932 7262 5944 7296
rect 5978 7262 5990 7296
rect 5932 7228 5990 7262
rect 5932 7194 5944 7228
rect 5978 7194 5990 7228
rect 5932 7160 5990 7194
rect 5932 7126 5944 7160
rect 5978 7126 5990 7160
rect 5932 7111 5990 7126
rect 6190 7296 6248 7311
rect 6190 7262 6202 7296
rect 6236 7262 6248 7296
rect 6190 7228 6248 7262
rect 6190 7194 6202 7228
rect 6236 7194 6248 7228
rect 6190 7160 6248 7194
rect 6190 7126 6202 7160
rect 6236 7126 6248 7160
rect 6190 7111 6248 7126
rect 3610 6878 3668 6893
rect 3610 6844 3622 6878
rect 3656 6844 3668 6878
rect 3610 6810 3668 6844
rect 3610 6776 3622 6810
rect 3656 6776 3668 6810
rect 3610 6742 3668 6776
rect 3610 6708 3622 6742
rect 3656 6708 3668 6742
rect 3610 6693 3668 6708
rect 3868 6878 3926 6893
rect 3868 6844 3880 6878
rect 3914 6844 3926 6878
rect 3868 6810 3926 6844
rect 3868 6776 3880 6810
rect 3914 6776 3926 6810
rect 3868 6742 3926 6776
rect 3868 6708 3880 6742
rect 3914 6708 3926 6742
rect 3868 6693 3926 6708
rect 4126 6878 4184 6893
rect 4126 6844 4138 6878
rect 4172 6844 4184 6878
rect 4126 6810 4184 6844
rect 4126 6776 4138 6810
rect 4172 6776 4184 6810
rect 4126 6742 4184 6776
rect 4126 6708 4138 6742
rect 4172 6708 4184 6742
rect 4126 6693 4184 6708
rect 4384 6878 4442 6893
rect 4384 6844 4396 6878
rect 4430 6844 4442 6878
rect 4384 6810 4442 6844
rect 4384 6776 4396 6810
rect 4430 6776 4442 6810
rect 4384 6742 4442 6776
rect 4384 6708 4396 6742
rect 4430 6708 4442 6742
rect 4384 6693 4442 6708
rect 4642 6878 4700 6893
rect 4642 6844 4654 6878
rect 4688 6844 4700 6878
rect 4642 6810 4700 6844
rect 4642 6776 4654 6810
rect 4688 6776 4700 6810
rect 4642 6742 4700 6776
rect 4642 6708 4654 6742
rect 4688 6708 4700 6742
rect 4642 6693 4700 6708
rect 4900 6878 4958 6893
rect 4900 6844 4912 6878
rect 4946 6844 4958 6878
rect 4900 6810 4958 6844
rect 4900 6776 4912 6810
rect 4946 6776 4958 6810
rect 4900 6742 4958 6776
rect 4900 6708 4912 6742
rect 4946 6708 4958 6742
rect 4900 6693 4958 6708
rect 5158 6878 5216 6893
rect 5158 6844 5170 6878
rect 5204 6844 5216 6878
rect 5158 6810 5216 6844
rect 5158 6776 5170 6810
rect 5204 6776 5216 6810
rect 5158 6742 5216 6776
rect 5158 6708 5170 6742
rect 5204 6708 5216 6742
rect 5158 6693 5216 6708
rect 5416 6878 5474 6893
rect 5416 6844 5428 6878
rect 5462 6844 5474 6878
rect 5416 6810 5474 6844
rect 5416 6776 5428 6810
rect 5462 6776 5474 6810
rect 5416 6742 5474 6776
rect 5416 6708 5428 6742
rect 5462 6708 5474 6742
rect 5416 6693 5474 6708
rect 5674 6878 5732 6893
rect 5674 6844 5686 6878
rect 5720 6844 5732 6878
rect 5674 6810 5732 6844
rect 5674 6776 5686 6810
rect 5720 6776 5732 6810
rect 5674 6742 5732 6776
rect 5674 6708 5686 6742
rect 5720 6708 5732 6742
rect 5674 6693 5732 6708
rect 5932 6878 5990 6893
rect 5932 6844 5944 6878
rect 5978 6844 5990 6878
rect 5932 6810 5990 6844
rect 5932 6776 5944 6810
rect 5978 6776 5990 6810
rect 5932 6742 5990 6776
rect 5932 6708 5944 6742
rect 5978 6708 5990 6742
rect 5932 6693 5990 6708
rect 6190 6878 6248 6893
rect 6190 6844 6202 6878
rect 6236 6844 6248 6878
rect 6190 6810 6248 6844
rect 6190 6776 6202 6810
rect 6236 6776 6248 6810
rect 6190 6742 6248 6776
rect 6190 6708 6202 6742
rect 6236 6708 6248 6742
rect 6190 6693 6248 6708
rect 3610 6460 3668 6475
rect 3610 6426 3622 6460
rect 3656 6426 3668 6460
rect 3610 6392 3668 6426
rect 3610 6358 3622 6392
rect 3656 6358 3668 6392
rect 3610 6324 3668 6358
rect 3610 6290 3622 6324
rect 3656 6290 3668 6324
rect 3610 6275 3668 6290
rect 3868 6460 3926 6475
rect 3868 6426 3880 6460
rect 3914 6426 3926 6460
rect 3868 6392 3926 6426
rect 3868 6358 3880 6392
rect 3914 6358 3926 6392
rect 3868 6324 3926 6358
rect 3868 6290 3880 6324
rect 3914 6290 3926 6324
rect 3868 6275 3926 6290
rect 4126 6460 4184 6475
rect 4126 6426 4138 6460
rect 4172 6426 4184 6460
rect 4126 6392 4184 6426
rect 4126 6358 4138 6392
rect 4172 6358 4184 6392
rect 4126 6324 4184 6358
rect 4126 6290 4138 6324
rect 4172 6290 4184 6324
rect 4126 6275 4184 6290
rect 4384 6460 4442 6475
rect 4384 6426 4396 6460
rect 4430 6426 4442 6460
rect 4384 6392 4442 6426
rect 4384 6358 4396 6392
rect 4430 6358 4442 6392
rect 4384 6324 4442 6358
rect 4384 6290 4396 6324
rect 4430 6290 4442 6324
rect 4384 6275 4442 6290
rect 4642 6460 4700 6475
rect 4642 6426 4654 6460
rect 4688 6426 4700 6460
rect 4642 6392 4700 6426
rect 4642 6358 4654 6392
rect 4688 6358 4700 6392
rect 4642 6324 4700 6358
rect 4642 6290 4654 6324
rect 4688 6290 4700 6324
rect 4642 6275 4700 6290
rect 4900 6460 4958 6475
rect 4900 6426 4912 6460
rect 4946 6426 4958 6460
rect 4900 6392 4958 6426
rect 4900 6358 4912 6392
rect 4946 6358 4958 6392
rect 4900 6324 4958 6358
rect 4900 6290 4912 6324
rect 4946 6290 4958 6324
rect 4900 6275 4958 6290
rect 5158 6460 5216 6475
rect 5158 6426 5170 6460
rect 5204 6426 5216 6460
rect 5158 6392 5216 6426
rect 5158 6358 5170 6392
rect 5204 6358 5216 6392
rect 5158 6324 5216 6358
rect 5158 6290 5170 6324
rect 5204 6290 5216 6324
rect 5158 6275 5216 6290
rect 5416 6460 5474 6475
rect 5416 6426 5428 6460
rect 5462 6426 5474 6460
rect 5416 6392 5474 6426
rect 5416 6358 5428 6392
rect 5462 6358 5474 6392
rect 5416 6324 5474 6358
rect 5416 6290 5428 6324
rect 5462 6290 5474 6324
rect 5416 6275 5474 6290
rect 5674 6460 5732 6475
rect 5674 6426 5686 6460
rect 5720 6426 5732 6460
rect 5674 6392 5732 6426
rect 5674 6358 5686 6392
rect 5720 6358 5732 6392
rect 5674 6324 5732 6358
rect 5674 6290 5686 6324
rect 5720 6290 5732 6324
rect 5674 6275 5732 6290
rect 5932 6460 5990 6475
rect 5932 6426 5944 6460
rect 5978 6426 5990 6460
rect 5932 6392 5990 6426
rect 5932 6358 5944 6392
rect 5978 6358 5990 6392
rect 5932 6324 5990 6358
rect 5932 6290 5944 6324
rect 5978 6290 5990 6324
rect 5932 6275 5990 6290
rect 6190 6460 6248 6475
rect 6190 6426 6202 6460
rect 6236 6426 6248 6460
rect 6190 6392 6248 6426
rect 6190 6358 6202 6392
rect 6236 6358 6248 6392
rect 6190 6324 6248 6358
rect 6190 6290 6202 6324
rect 6236 6290 6248 6324
rect 6190 6275 6248 6290
rect 3610 6042 3668 6057
rect 3610 6008 3622 6042
rect 3656 6008 3668 6042
rect 3610 5974 3668 6008
rect 3610 5940 3622 5974
rect 3656 5940 3668 5974
rect 3610 5906 3668 5940
rect 3610 5872 3622 5906
rect 3656 5872 3668 5906
rect 3610 5857 3668 5872
rect 3868 6042 3926 6057
rect 3868 6008 3880 6042
rect 3914 6008 3926 6042
rect 3868 5974 3926 6008
rect 3868 5940 3880 5974
rect 3914 5940 3926 5974
rect 3868 5906 3926 5940
rect 3868 5872 3880 5906
rect 3914 5872 3926 5906
rect 3868 5857 3926 5872
rect 4126 6042 4184 6057
rect 4126 6008 4138 6042
rect 4172 6008 4184 6042
rect 4126 5974 4184 6008
rect 4126 5940 4138 5974
rect 4172 5940 4184 5974
rect 4126 5906 4184 5940
rect 4126 5872 4138 5906
rect 4172 5872 4184 5906
rect 4126 5857 4184 5872
rect 4384 6042 4442 6057
rect 4384 6008 4396 6042
rect 4430 6008 4442 6042
rect 4384 5974 4442 6008
rect 4384 5940 4396 5974
rect 4430 5940 4442 5974
rect 4384 5906 4442 5940
rect 4384 5872 4396 5906
rect 4430 5872 4442 5906
rect 4384 5857 4442 5872
rect 4642 6042 4700 6057
rect 4642 6008 4654 6042
rect 4688 6008 4700 6042
rect 4642 5974 4700 6008
rect 4642 5940 4654 5974
rect 4688 5940 4700 5974
rect 4642 5906 4700 5940
rect 4642 5872 4654 5906
rect 4688 5872 4700 5906
rect 4642 5857 4700 5872
rect 4900 6042 4958 6057
rect 4900 6008 4912 6042
rect 4946 6008 4958 6042
rect 4900 5974 4958 6008
rect 4900 5940 4912 5974
rect 4946 5940 4958 5974
rect 4900 5906 4958 5940
rect 4900 5872 4912 5906
rect 4946 5872 4958 5906
rect 4900 5857 4958 5872
rect 5158 6042 5216 6057
rect 5158 6008 5170 6042
rect 5204 6008 5216 6042
rect 5158 5974 5216 6008
rect 5158 5940 5170 5974
rect 5204 5940 5216 5974
rect 5158 5906 5216 5940
rect 5158 5872 5170 5906
rect 5204 5872 5216 5906
rect 5158 5857 5216 5872
rect 5416 6042 5474 6057
rect 5416 6008 5428 6042
rect 5462 6008 5474 6042
rect 5416 5974 5474 6008
rect 5416 5940 5428 5974
rect 5462 5940 5474 5974
rect 5416 5906 5474 5940
rect 5416 5872 5428 5906
rect 5462 5872 5474 5906
rect 5416 5857 5474 5872
rect 5674 6042 5732 6057
rect 5674 6008 5686 6042
rect 5720 6008 5732 6042
rect 5674 5974 5732 6008
rect 5674 5940 5686 5974
rect 5720 5940 5732 5974
rect 5674 5906 5732 5940
rect 5674 5872 5686 5906
rect 5720 5872 5732 5906
rect 5674 5857 5732 5872
rect 5932 6042 5990 6057
rect 5932 6008 5944 6042
rect 5978 6008 5990 6042
rect 5932 5974 5990 6008
rect 5932 5940 5944 5974
rect 5978 5940 5990 5974
rect 5932 5906 5990 5940
rect 5932 5872 5944 5906
rect 5978 5872 5990 5906
rect 5932 5857 5990 5872
rect 6190 6042 6248 6057
rect 6190 6008 6202 6042
rect 6236 6008 6248 6042
rect 6190 5974 6248 6008
rect 6190 5940 6202 5974
rect 6236 5940 6248 5974
rect 6190 5906 6248 5940
rect 6190 5872 6202 5906
rect 6236 5872 6248 5906
rect 6190 5857 6248 5872
rect 3610 5624 3668 5639
rect 3610 5590 3622 5624
rect 3656 5590 3668 5624
rect 3610 5556 3668 5590
rect 3610 5522 3622 5556
rect 3656 5522 3668 5556
rect 3610 5488 3668 5522
rect 3610 5454 3622 5488
rect 3656 5454 3668 5488
rect 3610 5439 3668 5454
rect 3868 5624 3926 5639
rect 3868 5590 3880 5624
rect 3914 5590 3926 5624
rect 3868 5556 3926 5590
rect 3868 5522 3880 5556
rect 3914 5522 3926 5556
rect 3868 5488 3926 5522
rect 3868 5454 3880 5488
rect 3914 5454 3926 5488
rect 3868 5439 3926 5454
rect 4126 5624 4184 5639
rect 4126 5590 4138 5624
rect 4172 5590 4184 5624
rect 4126 5556 4184 5590
rect 4126 5522 4138 5556
rect 4172 5522 4184 5556
rect 4126 5488 4184 5522
rect 4126 5454 4138 5488
rect 4172 5454 4184 5488
rect 4126 5439 4184 5454
rect 4384 5624 4442 5639
rect 4384 5590 4396 5624
rect 4430 5590 4442 5624
rect 4384 5556 4442 5590
rect 4384 5522 4396 5556
rect 4430 5522 4442 5556
rect 4384 5488 4442 5522
rect 4384 5454 4396 5488
rect 4430 5454 4442 5488
rect 4384 5439 4442 5454
rect 4642 5624 4700 5639
rect 4642 5590 4654 5624
rect 4688 5590 4700 5624
rect 4642 5556 4700 5590
rect 4642 5522 4654 5556
rect 4688 5522 4700 5556
rect 4642 5488 4700 5522
rect 4642 5454 4654 5488
rect 4688 5454 4700 5488
rect 4642 5439 4700 5454
rect 4900 5624 4958 5639
rect 4900 5590 4912 5624
rect 4946 5590 4958 5624
rect 4900 5556 4958 5590
rect 4900 5522 4912 5556
rect 4946 5522 4958 5556
rect 4900 5488 4958 5522
rect 4900 5454 4912 5488
rect 4946 5454 4958 5488
rect 4900 5439 4958 5454
rect 5158 5624 5216 5639
rect 5158 5590 5170 5624
rect 5204 5590 5216 5624
rect 5158 5556 5216 5590
rect 5158 5522 5170 5556
rect 5204 5522 5216 5556
rect 5158 5488 5216 5522
rect 5158 5454 5170 5488
rect 5204 5454 5216 5488
rect 5158 5439 5216 5454
rect 5416 5624 5474 5639
rect 5416 5590 5428 5624
rect 5462 5590 5474 5624
rect 5416 5556 5474 5590
rect 5416 5522 5428 5556
rect 5462 5522 5474 5556
rect 5416 5488 5474 5522
rect 5416 5454 5428 5488
rect 5462 5454 5474 5488
rect 5416 5439 5474 5454
rect 5674 5624 5732 5639
rect 5674 5590 5686 5624
rect 5720 5590 5732 5624
rect 5674 5556 5732 5590
rect 5674 5522 5686 5556
rect 5720 5522 5732 5556
rect 5674 5488 5732 5522
rect 5674 5454 5686 5488
rect 5720 5454 5732 5488
rect 5674 5439 5732 5454
rect 5932 5624 5990 5639
rect 5932 5590 5944 5624
rect 5978 5590 5990 5624
rect 5932 5556 5990 5590
rect 5932 5522 5944 5556
rect 5978 5522 5990 5556
rect 5932 5488 5990 5522
rect 5932 5454 5944 5488
rect 5978 5454 5990 5488
rect 5932 5439 5990 5454
rect 6190 5624 6248 5639
rect 6190 5590 6202 5624
rect 6236 5590 6248 5624
rect 6190 5556 6248 5590
rect 6190 5522 6202 5556
rect 6236 5522 6248 5556
rect 6190 5488 6248 5522
rect 6190 5454 6202 5488
rect 6236 5454 6248 5488
rect 6190 5439 6248 5454
rect 3610 5206 3668 5221
rect 3610 5172 3622 5206
rect 3656 5172 3668 5206
rect 3610 5138 3668 5172
rect 3610 5104 3622 5138
rect 3656 5104 3668 5138
rect 3610 5070 3668 5104
rect 3610 5036 3622 5070
rect 3656 5036 3668 5070
rect 3610 5021 3668 5036
rect 3868 5206 3926 5221
rect 3868 5172 3880 5206
rect 3914 5172 3926 5206
rect 3868 5138 3926 5172
rect 3868 5104 3880 5138
rect 3914 5104 3926 5138
rect 3868 5070 3926 5104
rect 3868 5036 3880 5070
rect 3914 5036 3926 5070
rect 3868 5021 3926 5036
rect 4126 5206 4184 5221
rect 4126 5172 4138 5206
rect 4172 5172 4184 5206
rect 4126 5138 4184 5172
rect 4126 5104 4138 5138
rect 4172 5104 4184 5138
rect 4126 5070 4184 5104
rect 4126 5036 4138 5070
rect 4172 5036 4184 5070
rect 4126 5021 4184 5036
rect 4384 5206 4442 5221
rect 4384 5172 4396 5206
rect 4430 5172 4442 5206
rect 4384 5138 4442 5172
rect 4384 5104 4396 5138
rect 4430 5104 4442 5138
rect 4384 5070 4442 5104
rect 4384 5036 4396 5070
rect 4430 5036 4442 5070
rect 4384 5021 4442 5036
rect 4642 5206 4700 5221
rect 4642 5172 4654 5206
rect 4688 5172 4700 5206
rect 4642 5138 4700 5172
rect 4642 5104 4654 5138
rect 4688 5104 4700 5138
rect 4642 5070 4700 5104
rect 4642 5036 4654 5070
rect 4688 5036 4700 5070
rect 4642 5021 4700 5036
rect 4900 5206 4958 5221
rect 4900 5172 4912 5206
rect 4946 5172 4958 5206
rect 4900 5138 4958 5172
rect 4900 5104 4912 5138
rect 4946 5104 4958 5138
rect 4900 5070 4958 5104
rect 4900 5036 4912 5070
rect 4946 5036 4958 5070
rect 4900 5021 4958 5036
rect 5158 5206 5216 5221
rect 5158 5172 5170 5206
rect 5204 5172 5216 5206
rect 5158 5138 5216 5172
rect 5158 5104 5170 5138
rect 5204 5104 5216 5138
rect 5158 5070 5216 5104
rect 5158 5036 5170 5070
rect 5204 5036 5216 5070
rect 5158 5021 5216 5036
rect 5416 5206 5474 5221
rect 5416 5172 5428 5206
rect 5462 5172 5474 5206
rect 5416 5138 5474 5172
rect 5416 5104 5428 5138
rect 5462 5104 5474 5138
rect 5416 5070 5474 5104
rect 5416 5036 5428 5070
rect 5462 5036 5474 5070
rect 5416 5021 5474 5036
rect 5674 5206 5732 5221
rect 5674 5172 5686 5206
rect 5720 5172 5732 5206
rect 5674 5138 5732 5172
rect 5674 5104 5686 5138
rect 5720 5104 5732 5138
rect 5674 5070 5732 5104
rect 5674 5036 5686 5070
rect 5720 5036 5732 5070
rect 5674 5021 5732 5036
rect 5932 5206 5990 5221
rect 5932 5172 5944 5206
rect 5978 5172 5990 5206
rect 5932 5138 5990 5172
rect 5932 5104 5944 5138
rect 5978 5104 5990 5138
rect 5932 5070 5990 5104
rect 5932 5036 5944 5070
rect 5978 5036 5990 5070
rect 5932 5021 5990 5036
rect 6190 5206 6248 5221
rect 6190 5172 6202 5206
rect 6236 5172 6248 5206
rect 6190 5138 6248 5172
rect 6190 5104 6202 5138
rect 6236 5104 6248 5138
rect 6190 5070 6248 5104
rect 6190 5036 6202 5070
rect 6236 5036 6248 5070
rect 6190 5021 6248 5036
rect 3610 4788 3668 4803
rect 3610 4754 3622 4788
rect 3656 4754 3668 4788
rect 3610 4720 3668 4754
rect 3610 4686 3622 4720
rect 3656 4686 3668 4720
rect 3610 4652 3668 4686
rect 3610 4618 3622 4652
rect 3656 4618 3668 4652
rect 3610 4603 3668 4618
rect 3868 4788 3926 4803
rect 3868 4754 3880 4788
rect 3914 4754 3926 4788
rect 3868 4720 3926 4754
rect 3868 4686 3880 4720
rect 3914 4686 3926 4720
rect 3868 4652 3926 4686
rect 3868 4618 3880 4652
rect 3914 4618 3926 4652
rect 3868 4603 3926 4618
rect 4126 4788 4184 4803
rect 4126 4754 4138 4788
rect 4172 4754 4184 4788
rect 4126 4720 4184 4754
rect 4126 4686 4138 4720
rect 4172 4686 4184 4720
rect 4126 4652 4184 4686
rect 4126 4618 4138 4652
rect 4172 4618 4184 4652
rect 4126 4603 4184 4618
rect 4384 4788 4442 4803
rect 4384 4754 4396 4788
rect 4430 4754 4442 4788
rect 4384 4720 4442 4754
rect 4384 4686 4396 4720
rect 4430 4686 4442 4720
rect 4384 4652 4442 4686
rect 4384 4618 4396 4652
rect 4430 4618 4442 4652
rect 4384 4603 4442 4618
rect 4642 4788 4700 4803
rect 4642 4754 4654 4788
rect 4688 4754 4700 4788
rect 4642 4720 4700 4754
rect 4642 4686 4654 4720
rect 4688 4686 4700 4720
rect 4642 4652 4700 4686
rect 4642 4618 4654 4652
rect 4688 4618 4700 4652
rect 4642 4603 4700 4618
rect 4900 4788 4958 4803
rect 4900 4754 4912 4788
rect 4946 4754 4958 4788
rect 4900 4720 4958 4754
rect 4900 4686 4912 4720
rect 4946 4686 4958 4720
rect 4900 4652 4958 4686
rect 4900 4618 4912 4652
rect 4946 4618 4958 4652
rect 4900 4603 4958 4618
rect 5158 4788 5216 4803
rect 5158 4754 5170 4788
rect 5204 4754 5216 4788
rect 5158 4720 5216 4754
rect 5158 4686 5170 4720
rect 5204 4686 5216 4720
rect 5158 4652 5216 4686
rect 5158 4618 5170 4652
rect 5204 4618 5216 4652
rect 5158 4603 5216 4618
rect 5416 4788 5474 4803
rect 5416 4754 5428 4788
rect 5462 4754 5474 4788
rect 5416 4720 5474 4754
rect 5416 4686 5428 4720
rect 5462 4686 5474 4720
rect 5416 4652 5474 4686
rect 5416 4618 5428 4652
rect 5462 4618 5474 4652
rect 5416 4603 5474 4618
rect 5674 4788 5732 4803
rect 5674 4754 5686 4788
rect 5720 4754 5732 4788
rect 5674 4720 5732 4754
rect 5674 4686 5686 4720
rect 5720 4686 5732 4720
rect 5674 4652 5732 4686
rect 5674 4618 5686 4652
rect 5720 4618 5732 4652
rect 5674 4603 5732 4618
rect 5932 4788 5990 4803
rect 5932 4754 5944 4788
rect 5978 4754 5990 4788
rect 5932 4720 5990 4754
rect 5932 4686 5944 4720
rect 5978 4686 5990 4720
rect 5932 4652 5990 4686
rect 5932 4618 5944 4652
rect 5978 4618 5990 4652
rect 5932 4603 5990 4618
rect 6190 4788 6248 4803
rect 6190 4754 6202 4788
rect 6236 4754 6248 4788
rect 6190 4720 6248 4754
rect 6190 4686 6202 4720
rect 6236 4686 6248 4720
rect 6190 4652 6248 4686
rect 6190 4618 6202 4652
rect 6236 4618 6248 4652
rect 6190 4603 6248 4618
rect 3610 4370 3668 4385
rect 3610 4336 3622 4370
rect 3656 4336 3668 4370
rect 3610 4302 3668 4336
rect 3610 4268 3622 4302
rect 3656 4268 3668 4302
rect 3610 4234 3668 4268
rect 3610 4200 3622 4234
rect 3656 4200 3668 4234
rect 3610 4185 3668 4200
rect 3868 4370 3926 4385
rect 3868 4336 3880 4370
rect 3914 4336 3926 4370
rect 3868 4302 3926 4336
rect 3868 4268 3880 4302
rect 3914 4268 3926 4302
rect 3868 4234 3926 4268
rect 3868 4200 3880 4234
rect 3914 4200 3926 4234
rect 3868 4185 3926 4200
rect 4126 4370 4184 4385
rect 4126 4336 4138 4370
rect 4172 4336 4184 4370
rect 4126 4302 4184 4336
rect 4126 4268 4138 4302
rect 4172 4268 4184 4302
rect 4126 4234 4184 4268
rect 4126 4200 4138 4234
rect 4172 4200 4184 4234
rect 4126 4185 4184 4200
rect 4384 4370 4442 4385
rect 4384 4336 4396 4370
rect 4430 4336 4442 4370
rect 4384 4302 4442 4336
rect 4384 4268 4396 4302
rect 4430 4268 4442 4302
rect 4384 4234 4442 4268
rect 4384 4200 4396 4234
rect 4430 4200 4442 4234
rect 4384 4185 4442 4200
rect 4642 4370 4700 4385
rect 4642 4336 4654 4370
rect 4688 4336 4700 4370
rect 4642 4302 4700 4336
rect 4642 4268 4654 4302
rect 4688 4268 4700 4302
rect 4642 4234 4700 4268
rect 4642 4200 4654 4234
rect 4688 4200 4700 4234
rect 4642 4185 4700 4200
rect 4900 4370 4958 4385
rect 4900 4336 4912 4370
rect 4946 4336 4958 4370
rect 4900 4302 4958 4336
rect 4900 4268 4912 4302
rect 4946 4268 4958 4302
rect 4900 4234 4958 4268
rect 4900 4200 4912 4234
rect 4946 4200 4958 4234
rect 4900 4185 4958 4200
rect 5158 4370 5216 4385
rect 5158 4336 5170 4370
rect 5204 4336 5216 4370
rect 5158 4302 5216 4336
rect 5158 4268 5170 4302
rect 5204 4268 5216 4302
rect 5158 4234 5216 4268
rect 5158 4200 5170 4234
rect 5204 4200 5216 4234
rect 5158 4185 5216 4200
rect 5416 4370 5474 4385
rect 5416 4336 5428 4370
rect 5462 4336 5474 4370
rect 5416 4302 5474 4336
rect 5416 4268 5428 4302
rect 5462 4268 5474 4302
rect 5416 4234 5474 4268
rect 5416 4200 5428 4234
rect 5462 4200 5474 4234
rect 5416 4185 5474 4200
rect 5674 4370 5732 4385
rect 5674 4336 5686 4370
rect 5720 4336 5732 4370
rect 5674 4302 5732 4336
rect 5674 4268 5686 4302
rect 5720 4268 5732 4302
rect 5674 4234 5732 4268
rect 5674 4200 5686 4234
rect 5720 4200 5732 4234
rect 5674 4185 5732 4200
rect 5932 4370 5990 4385
rect 5932 4336 5944 4370
rect 5978 4336 5990 4370
rect 5932 4302 5990 4336
rect 5932 4268 5944 4302
rect 5978 4268 5990 4302
rect 5932 4234 5990 4268
rect 5932 4200 5944 4234
rect 5978 4200 5990 4234
rect 5932 4185 5990 4200
rect 6190 4370 6248 4385
rect 6190 4336 6202 4370
rect 6236 4336 6248 4370
rect 6190 4302 6248 4336
rect 6190 4268 6202 4302
rect 6236 4268 6248 4302
rect 6190 4234 6248 4268
rect 6190 4200 6202 4234
rect 6236 4200 6248 4234
rect 6190 4185 6248 4200
rect 8346 6885 8404 6900
rect 8346 6851 8358 6885
rect 8392 6851 8404 6885
rect 8346 6817 8404 6851
rect 8346 6783 8358 6817
rect 8392 6783 8404 6817
rect 8346 6749 8404 6783
rect 8346 6715 8358 6749
rect 8392 6715 8404 6749
rect 8346 6700 8404 6715
rect 8604 6885 8662 6900
rect 8604 6851 8616 6885
rect 8650 6851 8662 6885
rect 8604 6817 8662 6851
rect 8604 6783 8616 6817
rect 8650 6783 8662 6817
rect 8604 6749 8662 6783
rect 8604 6715 8616 6749
rect 8650 6715 8662 6749
rect 8604 6700 8662 6715
rect 8862 6885 8920 6900
rect 8862 6851 8874 6885
rect 8908 6851 8920 6885
rect 8862 6817 8920 6851
rect 8862 6783 8874 6817
rect 8908 6783 8920 6817
rect 8862 6749 8920 6783
rect 8862 6715 8874 6749
rect 8908 6715 8920 6749
rect 8862 6700 8920 6715
rect 9120 6885 9178 6900
rect 9120 6851 9132 6885
rect 9166 6851 9178 6885
rect 9120 6817 9178 6851
rect 9120 6783 9132 6817
rect 9166 6783 9178 6817
rect 9120 6749 9178 6783
rect 9120 6715 9132 6749
rect 9166 6715 9178 6749
rect 9120 6700 9178 6715
rect 9378 6885 9436 6900
rect 9378 6851 9390 6885
rect 9424 6851 9436 6885
rect 9378 6817 9436 6851
rect 9378 6783 9390 6817
rect 9424 6783 9436 6817
rect 9378 6749 9436 6783
rect 9378 6715 9390 6749
rect 9424 6715 9436 6749
rect 9378 6700 9436 6715
rect 9636 6885 9694 6900
rect 9636 6851 9648 6885
rect 9682 6851 9694 6885
rect 9636 6817 9694 6851
rect 9636 6783 9648 6817
rect 9682 6783 9694 6817
rect 9636 6749 9694 6783
rect 9636 6715 9648 6749
rect 9682 6715 9694 6749
rect 9636 6700 9694 6715
rect 9894 6885 9952 6900
rect 9894 6851 9906 6885
rect 9940 6851 9952 6885
rect 9894 6817 9952 6851
rect 9894 6783 9906 6817
rect 9940 6783 9952 6817
rect 9894 6749 9952 6783
rect 9894 6715 9906 6749
rect 9940 6715 9952 6749
rect 9894 6700 9952 6715
rect 8346 6467 8404 6482
rect 8346 6433 8358 6467
rect 8392 6433 8404 6467
rect 8346 6399 8404 6433
rect 8346 6365 8358 6399
rect 8392 6365 8404 6399
rect 8346 6331 8404 6365
rect 8346 6297 8358 6331
rect 8392 6297 8404 6331
rect 8346 6282 8404 6297
rect 8604 6467 8662 6482
rect 8604 6433 8616 6467
rect 8650 6433 8662 6467
rect 8604 6399 8662 6433
rect 8604 6365 8616 6399
rect 8650 6365 8662 6399
rect 8604 6331 8662 6365
rect 8604 6297 8616 6331
rect 8650 6297 8662 6331
rect 8604 6282 8662 6297
rect 8862 6467 8920 6482
rect 8862 6433 8874 6467
rect 8908 6433 8920 6467
rect 8862 6399 8920 6433
rect 8862 6365 8874 6399
rect 8908 6365 8920 6399
rect 8862 6331 8920 6365
rect 8862 6297 8874 6331
rect 8908 6297 8920 6331
rect 8862 6282 8920 6297
rect 9120 6467 9178 6482
rect 9120 6433 9132 6467
rect 9166 6433 9178 6467
rect 9120 6399 9178 6433
rect 9120 6365 9132 6399
rect 9166 6365 9178 6399
rect 9120 6331 9178 6365
rect 9120 6297 9132 6331
rect 9166 6297 9178 6331
rect 9120 6282 9178 6297
rect 9378 6467 9436 6482
rect 9378 6433 9390 6467
rect 9424 6433 9436 6467
rect 9378 6399 9436 6433
rect 9378 6365 9390 6399
rect 9424 6365 9436 6399
rect 9378 6331 9436 6365
rect 9378 6297 9390 6331
rect 9424 6297 9436 6331
rect 9378 6282 9436 6297
rect 9636 6467 9694 6482
rect 9636 6433 9648 6467
rect 9682 6433 9694 6467
rect 9636 6399 9694 6433
rect 9636 6365 9648 6399
rect 9682 6365 9694 6399
rect 9636 6331 9694 6365
rect 9636 6297 9648 6331
rect 9682 6297 9694 6331
rect 9636 6282 9694 6297
rect 9894 6467 9952 6482
rect 9894 6433 9906 6467
rect 9940 6433 9952 6467
rect 9894 6399 9952 6433
rect 9894 6365 9906 6399
rect 9940 6365 9952 6399
rect 9894 6331 9952 6365
rect 9894 6297 9906 6331
rect 9940 6297 9952 6331
rect 9894 6282 9952 6297
rect 8346 6049 8404 6064
rect 8346 6015 8358 6049
rect 8392 6015 8404 6049
rect 8346 5981 8404 6015
rect 8346 5947 8358 5981
rect 8392 5947 8404 5981
rect 8346 5913 8404 5947
rect 8346 5879 8358 5913
rect 8392 5879 8404 5913
rect 8346 5864 8404 5879
rect 8604 6049 8662 6064
rect 8604 6015 8616 6049
rect 8650 6015 8662 6049
rect 8604 5981 8662 6015
rect 8604 5947 8616 5981
rect 8650 5947 8662 5981
rect 8604 5913 8662 5947
rect 8604 5879 8616 5913
rect 8650 5879 8662 5913
rect 8604 5864 8662 5879
rect 8862 6049 8920 6064
rect 8862 6015 8874 6049
rect 8908 6015 8920 6049
rect 8862 5981 8920 6015
rect 8862 5947 8874 5981
rect 8908 5947 8920 5981
rect 8862 5913 8920 5947
rect 8862 5879 8874 5913
rect 8908 5879 8920 5913
rect 8862 5864 8920 5879
rect 9120 6049 9178 6064
rect 9120 6015 9132 6049
rect 9166 6015 9178 6049
rect 9120 5981 9178 6015
rect 9120 5947 9132 5981
rect 9166 5947 9178 5981
rect 9120 5913 9178 5947
rect 9120 5879 9132 5913
rect 9166 5879 9178 5913
rect 9120 5864 9178 5879
rect 9378 6049 9436 6064
rect 9378 6015 9390 6049
rect 9424 6015 9436 6049
rect 9378 5981 9436 6015
rect 9378 5947 9390 5981
rect 9424 5947 9436 5981
rect 9378 5913 9436 5947
rect 9378 5879 9390 5913
rect 9424 5879 9436 5913
rect 9378 5864 9436 5879
rect 9636 6049 9694 6064
rect 9636 6015 9648 6049
rect 9682 6015 9694 6049
rect 9636 5981 9694 6015
rect 9636 5947 9648 5981
rect 9682 5947 9694 5981
rect 9636 5913 9694 5947
rect 9636 5879 9648 5913
rect 9682 5879 9694 5913
rect 9636 5864 9694 5879
rect 9894 6049 9952 6064
rect 9894 6015 9906 6049
rect 9940 6015 9952 6049
rect 9894 5981 9952 6015
rect 9894 5947 9906 5981
rect 9940 5947 9952 5981
rect 9894 5913 9952 5947
rect 9894 5879 9906 5913
rect 9940 5879 9952 5913
rect 9894 5864 9952 5879
rect 8346 5631 8404 5646
rect 8346 5597 8358 5631
rect 8392 5597 8404 5631
rect 8346 5563 8404 5597
rect 8346 5529 8358 5563
rect 8392 5529 8404 5563
rect 8346 5495 8404 5529
rect 8346 5461 8358 5495
rect 8392 5461 8404 5495
rect 8346 5446 8404 5461
rect 8604 5631 8662 5646
rect 8604 5597 8616 5631
rect 8650 5597 8662 5631
rect 8604 5563 8662 5597
rect 8604 5529 8616 5563
rect 8650 5529 8662 5563
rect 8604 5495 8662 5529
rect 8604 5461 8616 5495
rect 8650 5461 8662 5495
rect 8604 5446 8662 5461
rect 8862 5631 8920 5646
rect 8862 5597 8874 5631
rect 8908 5597 8920 5631
rect 8862 5563 8920 5597
rect 8862 5529 8874 5563
rect 8908 5529 8920 5563
rect 8862 5495 8920 5529
rect 8862 5461 8874 5495
rect 8908 5461 8920 5495
rect 8862 5446 8920 5461
rect 9120 5631 9178 5646
rect 9120 5597 9132 5631
rect 9166 5597 9178 5631
rect 9120 5563 9178 5597
rect 9120 5529 9132 5563
rect 9166 5529 9178 5563
rect 9120 5495 9178 5529
rect 9120 5461 9132 5495
rect 9166 5461 9178 5495
rect 9120 5446 9178 5461
rect 9378 5631 9436 5646
rect 9378 5597 9390 5631
rect 9424 5597 9436 5631
rect 9378 5563 9436 5597
rect 9378 5529 9390 5563
rect 9424 5529 9436 5563
rect 9378 5495 9436 5529
rect 9378 5461 9390 5495
rect 9424 5461 9436 5495
rect 9378 5446 9436 5461
rect 9636 5631 9694 5646
rect 9636 5597 9648 5631
rect 9682 5597 9694 5631
rect 9636 5563 9694 5597
rect 9636 5529 9648 5563
rect 9682 5529 9694 5563
rect 9636 5495 9694 5529
rect 9636 5461 9648 5495
rect 9682 5461 9694 5495
rect 9636 5446 9694 5461
rect 9894 5631 9952 5646
rect 9894 5597 9906 5631
rect 9940 5597 9952 5631
rect 9894 5563 9952 5597
rect 9894 5529 9906 5563
rect 9940 5529 9952 5563
rect 9894 5495 9952 5529
rect 9894 5461 9906 5495
rect 9940 5461 9952 5495
rect 9894 5446 9952 5461
rect 8346 5213 8404 5228
rect 8346 5179 8358 5213
rect 8392 5179 8404 5213
rect 8346 5145 8404 5179
rect 8346 5111 8358 5145
rect 8392 5111 8404 5145
rect 8346 5077 8404 5111
rect 8346 5043 8358 5077
rect 8392 5043 8404 5077
rect 8346 5028 8404 5043
rect 8604 5213 8662 5228
rect 8604 5179 8616 5213
rect 8650 5179 8662 5213
rect 8604 5145 8662 5179
rect 8604 5111 8616 5145
rect 8650 5111 8662 5145
rect 8604 5077 8662 5111
rect 8604 5043 8616 5077
rect 8650 5043 8662 5077
rect 8604 5028 8662 5043
rect 8862 5213 8920 5228
rect 8862 5179 8874 5213
rect 8908 5179 8920 5213
rect 8862 5145 8920 5179
rect 8862 5111 8874 5145
rect 8908 5111 8920 5145
rect 8862 5077 8920 5111
rect 8862 5043 8874 5077
rect 8908 5043 8920 5077
rect 8862 5028 8920 5043
rect 9120 5213 9178 5228
rect 9120 5179 9132 5213
rect 9166 5179 9178 5213
rect 9120 5145 9178 5179
rect 9120 5111 9132 5145
rect 9166 5111 9178 5145
rect 9120 5077 9178 5111
rect 9120 5043 9132 5077
rect 9166 5043 9178 5077
rect 9120 5028 9178 5043
rect 9378 5213 9436 5228
rect 9378 5179 9390 5213
rect 9424 5179 9436 5213
rect 9378 5145 9436 5179
rect 9378 5111 9390 5145
rect 9424 5111 9436 5145
rect 9378 5077 9436 5111
rect 9378 5043 9390 5077
rect 9424 5043 9436 5077
rect 9378 5028 9436 5043
rect 9636 5213 9694 5228
rect 9636 5179 9648 5213
rect 9682 5179 9694 5213
rect 9636 5145 9694 5179
rect 9636 5111 9648 5145
rect 9682 5111 9694 5145
rect 9636 5077 9694 5111
rect 9636 5043 9648 5077
rect 9682 5043 9694 5077
rect 9636 5028 9694 5043
rect 9894 5213 9952 5228
rect 9894 5179 9906 5213
rect 9940 5179 9952 5213
rect 9894 5145 9952 5179
rect 9894 5111 9906 5145
rect 9940 5111 9952 5145
rect 9894 5077 9952 5111
rect 9894 5043 9906 5077
rect 9940 5043 9952 5077
rect 9894 5028 9952 5043
rect 8346 4795 8404 4810
rect 8346 4761 8358 4795
rect 8392 4761 8404 4795
rect 8346 4727 8404 4761
rect 8346 4693 8358 4727
rect 8392 4693 8404 4727
rect 8346 4659 8404 4693
rect 8346 4625 8358 4659
rect 8392 4625 8404 4659
rect 8346 4610 8404 4625
rect 8604 4795 8662 4810
rect 8604 4761 8616 4795
rect 8650 4761 8662 4795
rect 8604 4727 8662 4761
rect 8604 4693 8616 4727
rect 8650 4693 8662 4727
rect 8604 4659 8662 4693
rect 8604 4625 8616 4659
rect 8650 4625 8662 4659
rect 8604 4610 8662 4625
rect 8862 4795 8920 4810
rect 8862 4761 8874 4795
rect 8908 4761 8920 4795
rect 8862 4727 8920 4761
rect 8862 4693 8874 4727
rect 8908 4693 8920 4727
rect 8862 4659 8920 4693
rect 8862 4625 8874 4659
rect 8908 4625 8920 4659
rect 8862 4610 8920 4625
rect 9120 4795 9178 4810
rect 9120 4761 9132 4795
rect 9166 4761 9178 4795
rect 9120 4727 9178 4761
rect 9120 4693 9132 4727
rect 9166 4693 9178 4727
rect 9120 4659 9178 4693
rect 9120 4625 9132 4659
rect 9166 4625 9178 4659
rect 9120 4610 9178 4625
rect 9378 4795 9436 4810
rect 9378 4761 9390 4795
rect 9424 4761 9436 4795
rect 9378 4727 9436 4761
rect 9378 4693 9390 4727
rect 9424 4693 9436 4727
rect 9378 4659 9436 4693
rect 9378 4625 9390 4659
rect 9424 4625 9436 4659
rect 9378 4610 9436 4625
rect 9636 4795 9694 4810
rect 9636 4761 9648 4795
rect 9682 4761 9694 4795
rect 9636 4727 9694 4761
rect 9636 4693 9648 4727
rect 9682 4693 9694 4727
rect 9636 4659 9694 4693
rect 9636 4625 9648 4659
rect 9682 4625 9694 4659
rect 9636 4610 9694 4625
rect 9894 4795 9952 4810
rect 9894 4761 9906 4795
rect 9940 4761 9952 4795
rect 9894 4727 9952 4761
rect 9894 4693 9906 4727
rect 9940 4693 9952 4727
rect 9894 4659 9952 4693
rect 9894 4625 9906 4659
rect 9940 4625 9952 4659
rect 9894 4610 9952 4625
rect 8346 4377 8404 4392
rect 8346 4343 8358 4377
rect 8392 4343 8404 4377
rect 8346 4309 8404 4343
rect 8346 4275 8358 4309
rect 8392 4275 8404 4309
rect 8346 4241 8404 4275
rect 8346 4207 8358 4241
rect 8392 4207 8404 4241
rect 8346 4192 8404 4207
rect 8604 4377 8662 4392
rect 8604 4343 8616 4377
rect 8650 4343 8662 4377
rect 8604 4309 8662 4343
rect 8604 4275 8616 4309
rect 8650 4275 8662 4309
rect 8604 4241 8662 4275
rect 8604 4207 8616 4241
rect 8650 4207 8662 4241
rect 8604 4192 8662 4207
rect 8862 4377 8920 4392
rect 8862 4343 8874 4377
rect 8908 4343 8920 4377
rect 8862 4309 8920 4343
rect 8862 4275 8874 4309
rect 8908 4275 8920 4309
rect 8862 4241 8920 4275
rect 8862 4207 8874 4241
rect 8908 4207 8920 4241
rect 8862 4192 8920 4207
rect 9120 4377 9178 4392
rect 9120 4343 9132 4377
rect 9166 4343 9178 4377
rect 9120 4309 9178 4343
rect 9120 4275 9132 4309
rect 9166 4275 9178 4309
rect 9120 4241 9178 4275
rect 9120 4207 9132 4241
rect 9166 4207 9178 4241
rect 9120 4192 9178 4207
rect 9378 4377 9436 4392
rect 9378 4343 9390 4377
rect 9424 4343 9436 4377
rect 9378 4309 9436 4343
rect 9378 4275 9390 4309
rect 9424 4275 9436 4309
rect 9378 4241 9436 4275
rect 9378 4207 9390 4241
rect 9424 4207 9436 4241
rect 9378 4192 9436 4207
rect 9636 4377 9694 4392
rect 9636 4343 9648 4377
rect 9682 4343 9694 4377
rect 9636 4309 9694 4343
rect 9636 4275 9648 4309
rect 9682 4275 9694 4309
rect 9636 4241 9694 4275
rect 9636 4207 9648 4241
rect 9682 4207 9694 4241
rect 9636 4192 9694 4207
rect 9894 4377 9952 4392
rect 9894 4343 9906 4377
rect 9940 4343 9952 4377
rect 9894 4309 9952 4343
rect 9894 4275 9906 4309
rect 9940 4275 9952 4309
rect 9894 4241 9952 4275
rect 9894 4207 9906 4241
rect 9940 4207 9952 4241
rect 9894 4192 9952 4207
<< pdiff >>
rect -1251 10465 -1193 10480
rect -1251 10431 -1239 10465
rect -1205 10431 -1193 10465
rect -1251 10397 -1193 10431
rect -1251 10363 -1239 10397
rect -1205 10363 -1193 10397
rect -1251 10329 -1193 10363
rect -1251 10295 -1239 10329
rect -1205 10295 -1193 10329
rect -1251 10280 -1193 10295
rect -993 10465 -935 10480
rect -993 10431 -981 10465
rect -947 10431 -935 10465
rect -993 10397 -935 10431
rect -993 10363 -981 10397
rect -947 10363 -935 10397
rect -993 10329 -935 10363
rect -993 10295 -981 10329
rect -947 10295 -935 10329
rect -993 10280 -935 10295
rect -735 10465 -677 10480
rect -735 10431 -723 10465
rect -689 10431 -677 10465
rect -735 10397 -677 10431
rect -735 10363 -723 10397
rect -689 10363 -677 10397
rect -735 10329 -677 10363
rect -735 10295 -723 10329
rect -689 10295 -677 10329
rect -735 10280 -677 10295
rect -477 10465 -419 10480
rect -477 10431 -465 10465
rect -431 10431 -419 10465
rect -477 10397 -419 10431
rect -477 10363 -465 10397
rect -431 10363 -419 10397
rect -477 10329 -419 10363
rect -477 10295 -465 10329
rect -431 10295 -419 10329
rect -477 10280 -419 10295
rect -219 10465 -161 10480
rect -219 10431 -207 10465
rect -173 10431 -161 10465
rect -219 10397 -161 10431
rect -219 10363 -207 10397
rect -173 10363 -161 10397
rect -219 10329 -161 10363
rect -219 10295 -207 10329
rect -173 10295 -161 10329
rect -219 10280 -161 10295
rect 39 10465 97 10480
rect 39 10431 51 10465
rect 85 10431 97 10465
rect 39 10397 97 10431
rect 39 10363 51 10397
rect 85 10363 97 10397
rect 39 10329 97 10363
rect 39 10295 51 10329
rect 85 10295 97 10329
rect 39 10280 97 10295
rect 297 10465 355 10480
rect 297 10431 309 10465
rect 343 10431 355 10465
rect 297 10397 355 10431
rect 297 10363 309 10397
rect 343 10363 355 10397
rect 297 10329 355 10363
rect 297 10295 309 10329
rect 343 10295 355 10329
rect 297 10280 355 10295
rect -1251 10029 -1193 10044
rect -1251 9995 -1239 10029
rect -1205 9995 -1193 10029
rect -1251 9961 -1193 9995
rect -1251 9927 -1239 9961
rect -1205 9927 -1193 9961
rect -1251 9893 -1193 9927
rect -1251 9859 -1239 9893
rect -1205 9859 -1193 9893
rect -1251 9844 -1193 9859
rect -993 10029 -935 10044
rect -993 9995 -981 10029
rect -947 9995 -935 10029
rect -993 9961 -935 9995
rect -993 9927 -981 9961
rect -947 9927 -935 9961
rect -993 9893 -935 9927
rect -993 9859 -981 9893
rect -947 9859 -935 9893
rect -993 9844 -935 9859
rect -735 10029 -677 10044
rect -735 9995 -723 10029
rect -689 9995 -677 10029
rect -735 9961 -677 9995
rect -735 9927 -723 9961
rect -689 9927 -677 9961
rect -735 9893 -677 9927
rect -735 9859 -723 9893
rect -689 9859 -677 9893
rect -735 9844 -677 9859
rect -477 10029 -419 10044
rect -477 9995 -465 10029
rect -431 9995 -419 10029
rect -477 9961 -419 9995
rect -477 9927 -465 9961
rect -431 9927 -419 9961
rect -477 9893 -419 9927
rect -477 9859 -465 9893
rect -431 9859 -419 9893
rect -477 9844 -419 9859
rect -219 10029 -161 10044
rect -219 9995 -207 10029
rect -173 9995 -161 10029
rect -219 9961 -161 9995
rect -219 9927 -207 9961
rect -173 9927 -161 9961
rect -219 9893 -161 9927
rect -219 9859 -207 9893
rect -173 9859 -161 9893
rect -219 9844 -161 9859
rect 39 10029 97 10044
rect 39 9995 51 10029
rect 85 9995 97 10029
rect 39 9961 97 9995
rect 39 9927 51 9961
rect 85 9927 97 9961
rect 39 9893 97 9927
rect 39 9859 51 9893
rect 85 9859 97 9893
rect 39 9844 97 9859
rect 297 10029 355 10044
rect 297 9995 309 10029
rect 343 9995 355 10029
rect 297 9961 355 9995
rect 297 9927 309 9961
rect 343 9927 355 9961
rect 297 9893 355 9927
rect 297 9859 309 9893
rect 343 9859 355 9893
rect 297 9844 355 9859
rect -1251 9593 -1193 9608
rect -1251 9559 -1239 9593
rect -1205 9559 -1193 9593
rect -1251 9525 -1193 9559
rect -1251 9491 -1239 9525
rect -1205 9491 -1193 9525
rect -1251 9457 -1193 9491
rect -1251 9423 -1239 9457
rect -1205 9423 -1193 9457
rect -1251 9408 -1193 9423
rect -993 9593 -935 9608
rect -993 9559 -981 9593
rect -947 9559 -935 9593
rect -993 9525 -935 9559
rect -993 9491 -981 9525
rect -947 9491 -935 9525
rect -993 9457 -935 9491
rect -993 9423 -981 9457
rect -947 9423 -935 9457
rect -993 9408 -935 9423
rect -735 9593 -677 9608
rect -735 9559 -723 9593
rect -689 9559 -677 9593
rect -735 9525 -677 9559
rect -735 9491 -723 9525
rect -689 9491 -677 9525
rect -735 9457 -677 9491
rect -735 9423 -723 9457
rect -689 9423 -677 9457
rect -735 9408 -677 9423
rect -477 9593 -419 9608
rect -477 9559 -465 9593
rect -431 9559 -419 9593
rect -477 9525 -419 9559
rect -477 9491 -465 9525
rect -431 9491 -419 9525
rect -477 9457 -419 9491
rect -477 9423 -465 9457
rect -431 9423 -419 9457
rect -477 9408 -419 9423
rect -219 9593 -161 9608
rect -219 9559 -207 9593
rect -173 9559 -161 9593
rect -219 9525 -161 9559
rect -219 9491 -207 9525
rect -173 9491 -161 9525
rect -219 9457 -161 9491
rect -219 9423 -207 9457
rect -173 9423 -161 9457
rect -219 9408 -161 9423
rect 39 9593 97 9608
rect 39 9559 51 9593
rect 85 9559 97 9593
rect 39 9525 97 9559
rect 39 9491 51 9525
rect 85 9491 97 9525
rect 39 9457 97 9491
rect 39 9423 51 9457
rect 85 9423 97 9457
rect 39 9408 97 9423
rect 297 9593 355 9608
rect 297 9559 309 9593
rect 343 9559 355 9593
rect 297 9525 355 9559
rect 297 9491 309 9525
rect 343 9491 355 9525
rect 297 9457 355 9491
rect 297 9423 309 9457
rect 343 9423 355 9457
rect 297 9408 355 9423
rect -1251 9157 -1193 9172
rect -1251 9123 -1239 9157
rect -1205 9123 -1193 9157
rect -1251 9089 -1193 9123
rect -1251 9055 -1239 9089
rect -1205 9055 -1193 9089
rect -1251 9021 -1193 9055
rect -1251 8987 -1239 9021
rect -1205 8987 -1193 9021
rect -1251 8972 -1193 8987
rect -993 9157 -935 9172
rect -993 9123 -981 9157
rect -947 9123 -935 9157
rect -993 9089 -935 9123
rect -993 9055 -981 9089
rect -947 9055 -935 9089
rect -993 9021 -935 9055
rect -993 8987 -981 9021
rect -947 8987 -935 9021
rect -993 8972 -935 8987
rect -735 9157 -677 9172
rect -735 9123 -723 9157
rect -689 9123 -677 9157
rect -735 9089 -677 9123
rect -735 9055 -723 9089
rect -689 9055 -677 9089
rect -735 9021 -677 9055
rect -735 8987 -723 9021
rect -689 8987 -677 9021
rect -735 8972 -677 8987
rect -477 9157 -419 9172
rect -477 9123 -465 9157
rect -431 9123 -419 9157
rect -477 9089 -419 9123
rect -477 9055 -465 9089
rect -431 9055 -419 9089
rect -477 9021 -419 9055
rect -477 8987 -465 9021
rect -431 8987 -419 9021
rect -477 8972 -419 8987
rect -219 9157 -161 9172
rect -219 9123 -207 9157
rect -173 9123 -161 9157
rect -219 9089 -161 9123
rect -219 9055 -207 9089
rect -173 9055 -161 9089
rect -219 9021 -161 9055
rect -219 8987 -207 9021
rect -173 8987 -161 9021
rect -219 8972 -161 8987
rect 39 9157 97 9172
rect 39 9123 51 9157
rect 85 9123 97 9157
rect 39 9089 97 9123
rect 39 9055 51 9089
rect 85 9055 97 9089
rect 39 9021 97 9055
rect 39 8987 51 9021
rect 85 8987 97 9021
rect 39 8972 97 8987
rect 297 9157 355 9172
rect 297 9123 309 9157
rect 343 9123 355 9157
rect 297 9089 355 9123
rect 297 9055 309 9089
rect 343 9055 355 9089
rect 297 9021 355 9055
rect 297 8987 309 9021
rect 343 8987 355 9021
rect 297 8972 355 8987
rect 6997 10783 7055 10798
rect 6997 10749 7009 10783
rect 7043 10749 7055 10783
rect 6997 10715 7055 10749
rect 6997 10681 7009 10715
rect 7043 10681 7055 10715
rect 6997 10647 7055 10681
rect 6997 10613 7009 10647
rect 7043 10613 7055 10647
rect 6997 10598 7055 10613
rect 7255 10783 7313 10798
rect 7255 10749 7267 10783
rect 7301 10749 7313 10783
rect 7255 10715 7313 10749
rect 7255 10681 7267 10715
rect 7301 10681 7313 10715
rect 7255 10647 7313 10681
rect 7255 10613 7267 10647
rect 7301 10613 7313 10647
rect 7255 10598 7313 10613
rect 7513 10783 7571 10798
rect 7513 10749 7525 10783
rect 7559 10749 7571 10783
rect 7513 10715 7571 10749
rect 7513 10681 7525 10715
rect 7559 10681 7571 10715
rect 7513 10647 7571 10681
rect 7513 10613 7525 10647
rect 7559 10613 7571 10647
rect 7513 10598 7571 10613
rect 7771 10783 7829 10798
rect 7771 10749 7783 10783
rect 7817 10749 7829 10783
rect 7771 10715 7829 10749
rect 7771 10681 7783 10715
rect 7817 10681 7829 10715
rect 7771 10647 7829 10681
rect 7771 10613 7783 10647
rect 7817 10613 7829 10647
rect 7771 10598 7829 10613
rect 8029 10783 8087 10798
rect 8029 10749 8041 10783
rect 8075 10749 8087 10783
rect 8029 10715 8087 10749
rect 8029 10681 8041 10715
rect 8075 10681 8087 10715
rect 8029 10647 8087 10681
rect 8029 10613 8041 10647
rect 8075 10613 8087 10647
rect 8029 10598 8087 10613
rect 8287 10783 8345 10798
rect 8287 10749 8299 10783
rect 8333 10749 8345 10783
rect 8287 10715 8345 10749
rect 8287 10681 8299 10715
rect 8333 10681 8345 10715
rect 8287 10647 8345 10681
rect 8287 10613 8299 10647
rect 8333 10613 8345 10647
rect 8287 10598 8345 10613
rect 8545 10783 8603 10798
rect 8545 10749 8557 10783
rect 8591 10749 8603 10783
rect 8545 10715 8603 10749
rect 8545 10681 8557 10715
rect 8591 10681 8603 10715
rect 8545 10647 8603 10681
rect 8545 10613 8557 10647
rect 8591 10613 8603 10647
rect 8545 10598 8603 10613
rect 6997 10347 7055 10362
rect 6997 10313 7009 10347
rect 7043 10313 7055 10347
rect 6997 10279 7055 10313
rect 6997 10245 7009 10279
rect 7043 10245 7055 10279
rect 6997 10211 7055 10245
rect 6997 10177 7009 10211
rect 7043 10177 7055 10211
rect 6997 10162 7055 10177
rect 7255 10347 7313 10362
rect 7255 10313 7267 10347
rect 7301 10313 7313 10347
rect 7255 10279 7313 10313
rect 7255 10245 7267 10279
rect 7301 10245 7313 10279
rect 7255 10211 7313 10245
rect 7255 10177 7267 10211
rect 7301 10177 7313 10211
rect 7255 10162 7313 10177
rect 7513 10347 7571 10362
rect 7513 10313 7525 10347
rect 7559 10313 7571 10347
rect 7513 10279 7571 10313
rect 7513 10245 7525 10279
rect 7559 10245 7571 10279
rect 7513 10211 7571 10245
rect 7513 10177 7525 10211
rect 7559 10177 7571 10211
rect 7513 10162 7571 10177
rect 7771 10347 7829 10362
rect 7771 10313 7783 10347
rect 7817 10313 7829 10347
rect 7771 10279 7829 10313
rect 7771 10245 7783 10279
rect 7817 10245 7829 10279
rect 7771 10211 7829 10245
rect 7771 10177 7783 10211
rect 7817 10177 7829 10211
rect 7771 10162 7829 10177
rect 8029 10347 8087 10362
rect 8029 10313 8041 10347
rect 8075 10313 8087 10347
rect 8029 10279 8087 10313
rect 8029 10245 8041 10279
rect 8075 10245 8087 10279
rect 8029 10211 8087 10245
rect 8029 10177 8041 10211
rect 8075 10177 8087 10211
rect 8029 10162 8087 10177
rect 8287 10347 8345 10362
rect 8287 10313 8299 10347
rect 8333 10313 8345 10347
rect 8287 10279 8345 10313
rect 8287 10245 8299 10279
rect 8333 10245 8345 10279
rect 8287 10211 8345 10245
rect 8287 10177 8299 10211
rect 8333 10177 8345 10211
rect 8287 10162 8345 10177
rect 8545 10347 8603 10362
rect 8545 10313 8557 10347
rect 8591 10313 8603 10347
rect 8545 10279 8603 10313
rect 8545 10245 8557 10279
rect 8591 10245 8603 10279
rect 8545 10211 8603 10245
rect 8545 10177 8557 10211
rect 8591 10177 8603 10211
rect 8545 10162 8603 10177
rect 6997 9911 7055 9926
rect 6997 9877 7009 9911
rect 7043 9877 7055 9911
rect 6997 9843 7055 9877
rect 6997 9809 7009 9843
rect 7043 9809 7055 9843
rect 6997 9775 7055 9809
rect 6997 9741 7009 9775
rect 7043 9741 7055 9775
rect 6997 9726 7055 9741
rect 7255 9911 7313 9926
rect 7255 9877 7267 9911
rect 7301 9877 7313 9911
rect 7255 9843 7313 9877
rect 7255 9809 7267 9843
rect 7301 9809 7313 9843
rect 7255 9775 7313 9809
rect 7255 9741 7267 9775
rect 7301 9741 7313 9775
rect 7255 9726 7313 9741
rect 7513 9911 7571 9926
rect 7513 9877 7525 9911
rect 7559 9877 7571 9911
rect 7513 9843 7571 9877
rect 7513 9809 7525 9843
rect 7559 9809 7571 9843
rect 7513 9775 7571 9809
rect 7513 9741 7525 9775
rect 7559 9741 7571 9775
rect 7513 9726 7571 9741
rect 7771 9911 7829 9926
rect 7771 9877 7783 9911
rect 7817 9877 7829 9911
rect 7771 9843 7829 9877
rect 7771 9809 7783 9843
rect 7817 9809 7829 9843
rect 7771 9775 7829 9809
rect 7771 9741 7783 9775
rect 7817 9741 7829 9775
rect 7771 9726 7829 9741
rect 8029 9911 8087 9926
rect 8029 9877 8041 9911
rect 8075 9877 8087 9911
rect 8029 9843 8087 9877
rect 8029 9809 8041 9843
rect 8075 9809 8087 9843
rect 8029 9775 8087 9809
rect 8029 9741 8041 9775
rect 8075 9741 8087 9775
rect 8029 9726 8087 9741
rect 8287 9911 8345 9926
rect 8287 9877 8299 9911
rect 8333 9877 8345 9911
rect 8287 9843 8345 9877
rect 8287 9809 8299 9843
rect 8333 9809 8345 9843
rect 8287 9775 8345 9809
rect 8287 9741 8299 9775
rect 8333 9741 8345 9775
rect 8287 9726 8345 9741
rect 8545 9911 8603 9926
rect 8545 9877 8557 9911
rect 8591 9877 8603 9911
rect 8545 9843 8603 9877
rect 8545 9809 8557 9843
rect 8591 9809 8603 9843
rect 8545 9775 8603 9809
rect 8545 9741 8557 9775
rect 8591 9741 8603 9775
rect 8545 9726 8603 9741
rect 6997 9475 7055 9490
rect 6997 9441 7009 9475
rect 7043 9441 7055 9475
rect 6997 9407 7055 9441
rect 6997 9373 7009 9407
rect 7043 9373 7055 9407
rect 6997 9339 7055 9373
rect 6997 9305 7009 9339
rect 7043 9305 7055 9339
rect 6997 9290 7055 9305
rect 7255 9475 7313 9490
rect 7255 9441 7267 9475
rect 7301 9441 7313 9475
rect 7255 9407 7313 9441
rect 7255 9373 7267 9407
rect 7301 9373 7313 9407
rect 7255 9339 7313 9373
rect 7255 9305 7267 9339
rect 7301 9305 7313 9339
rect 7255 9290 7313 9305
rect 7513 9475 7571 9490
rect 7513 9441 7525 9475
rect 7559 9441 7571 9475
rect 7513 9407 7571 9441
rect 7513 9373 7525 9407
rect 7559 9373 7571 9407
rect 7513 9339 7571 9373
rect 7513 9305 7525 9339
rect 7559 9305 7571 9339
rect 7513 9290 7571 9305
rect 7771 9475 7829 9490
rect 7771 9441 7783 9475
rect 7817 9441 7829 9475
rect 7771 9407 7829 9441
rect 7771 9373 7783 9407
rect 7817 9373 7829 9407
rect 7771 9339 7829 9373
rect 7771 9305 7783 9339
rect 7817 9305 7829 9339
rect 7771 9290 7829 9305
rect 8029 9475 8087 9490
rect 8029 9441 8041 9475
rect 8075 9441 8087 9475
rect 8029 9407 8087 9441
rect 8029 9373 8041 9407
rect 8075 9373 8087 9407
rect 8029 9339 8087 9373
rect 8029 9305 8041 9339
rect 8075 9305 8087 9339
rect 8029 9290 8087 9305
rect 8287 9475 8345 9490
rect 8287 9441 8299 9475
rect 8333 9441 8345 9475
rect 8287 9407 8345 9441
rect 8287 9373 8299 9407
rect 8333 9373 8345 9407
rect 8287 9339 8345 9373
rect 8287 9305 8299 9339
rect 8333 9305 8345 9339
rect 8287 9290 8345 9305
rect 8545 9475 8603 9490
rect 8545 9441 8557 9475
rect 8591 9441 8603 9475
rect 8545 9407 8603 9441
rect 8545 9373 8557 9407
rect 8591 9373 8603 9407
rect 8545 9339 8603 9373
rect 8545 9305 8557 9339
rect 8591 9305 8603 9339
rect 8545 9290 8603 9305
rect 6997 9039 7055 9054
rect 6997 9005 7009 9039
rect 7043 9005 7055 9039
rect 6997 8971 7055 9005
rect 6997 8937 7009 8971
rect 7043 8937 7055 8971
rect 6997 8903 7055 8937
rect 6997 8869 7009 8903
rect 7043 8869 7055 8903
rect 6997 8854 7055 8869
rect 7255 9039 7313 9054
rect 7255 9005 7267 9039
rect 7301 9005 7313 9039
rect 7255 8971 7313 9005
rect 7255 8937 7267 8971
rect 7301 8937 7313 8971
rect 7255 8903 7313 8937
rect 7255 8869 7267 8903
rect 7301 8869 7313 8903
rect 7255 8854 7313 8869
rect 7513 9039 7571 9054
rect 7513 9005 7525 9039
rect 7559 9005 7571 9039
rect 7513 8971 7571 9005
rect 7513 8937 7525 8971
rect 7559 8937 7571 8971
rect 7513 8903 7571 8937
rect 7513 8869 7525 8903
rect 7559 8869 7571 8903
rect 7513 8854 7571 8869
rect 7771 9039 7829 9054
rect 7771 9005 7783 9039
rect 7817 9005 7829 9039
rect 7771 8971 7829 9005
rect 7771 8937 7783 8971
rect 7817 8937 7829 8971
rect 7771 8903 7829 8937
rect 7771 8869 7783 8903
rect 7817 8869 7829 8903
rect 7771 8854 7829 8869
rect 8029 9039 8087 9054
rect 8029 9005 8041 9039
rect 8075 9005 8087 9039
rect 8029 8971 8087 9005
rect 8029 8937 8041 8971
rect 8075 8937 8087 8971
rect 8029 8903 8087 8937
rect 8029 8869 8041 8903
rect 8075 8869 8087 8903
rect 8029 8854 8087 8869
rect 8287 9039 8345 9054
rect 8287 9005 8299 9039
rect 8333 9005 8345 9039
rect 8287 8971 8345 9005
rect 8287 8937 8299 8971
rect 8333 8937 8345 8971
rect 8287 8903 8345 8937
rect 8287 8869 8299 8903
rect 8333 8869 8345 8903
rect 8287 8854 8345 8869
rect 8545 9039 8603 9054
rect 8545 9005 8557 9039
rect 8591 9005 8603 9039
rect 8545 8971 8603 9005
rect 8545 8937 8557 8971
rect 8591 8937 8603 8971
rect 8545 8903 8603 8937
rect 8545 8869 8557 8903
rect 8591 8869 8603 8903
rect 8545 8854 8603 8869
rect 6997 8603 7055 8618
rect 6997 8569 7009 8603
rect 7043 8569 7055 8603
rect 6997 8535 7055 8569
rect 6997 8501 7009 8535
rect 7043 8501 7055 8535
rect 6997 8467 7055 8501
rect 6997 8433 7009 8467
rect 7043 8433 7055 8467
rect 6997 8418 7055 8433
rect 7255 8603 7313 8618
rect 7255 8569 7267 8603
rect 7301 8569 7313 8603
rect 7255 8535 7313 8569
rect 7255 8501 7267 8535
rect 7301 8501 7313 8535
rect 7255 8467 7313 8501
rect 7255 8433 7267 8467
rect 7301 8433 7313 8467
rect 7255 8418 7313 8433
rect 7513 8603 7571 8618
rect 7513 8569 7525 8603
rect 7559 8569 7571 8603
rect 7513 8535 7571 8569
rect 7513 8501 7525 8535
rect 7559 8501 7571 8535
rect 7513 8467 7571 8501
rect 7513 8433 7525 8467
rect 7559 8433 7571 8467
rect 7513 8418 7571 8433
rect 7771 8603 7829 8618
rect 7771 8569 7783 8603
rect 7817 8569 7829 8603
rect 7771 8535 7829 8569
rect 7771 8501 7783 8535
rect 7817 8501 7829 8535
rect 7771 8467 7829 8501
rect 7771 8433 7783 8467
rect 7817 8433 7829 8467
rect 7771 8418 7829 8433
rect 8029 8603 8087 8618
rect 8029 8569 8041 8603
rect 8075 8569 8087 8603
rect 8029 8535 8087 8569
rect 8029 8501 8041 8535
rect 8075 8501 8087 8535
rect 8029 8467 8087 8501
rect 8029 8433 8041 8467
rect 8075 8433 8087 8467
rect 8029 8418 8087 8433
rect 8287 8603 8345 8618
rect 8287 8569 8299 8603
rect 8333 8569 8345 8603
rect 8287 8535 8345 8569
rect 8287 8501 8299 8535
rect 8333 8501 8345 8535
rect 8287 8467 8345 8501
rect 8287 8433 8299 8467
rect 8333 8433 8345 8467
rect 8287 8418 8345 8433
rect 8545 8603 8603 8618
rect 8545 8569 8557 8603
rect 8591 8569 8603 8603
rect 8545 8535 8603 8569
rect 8545 8501 8557 8535
rect 8591 8501 8603 8535
rect 8545 8467 8603 8501
rect 8545 8433 8557 8467
rect 8591 8433 8603 8467
rect 8545 8418 8603 8433
rect 6997 8167 7055 8182
rect 6997 8133 7009 8167
rect 7043 8133 7055 8167
rect 6997 8099 7055 8133
rect 6997 8065 7009 8099
rect 7043 8065 7055 8099
rect 6997 8031 7055 8065
rect 6997 7997 7009 8031
rect 7043 7997 7055 8031
rect 6997 7982 7055 7997
rect 7255 8167 7313 8182
rect 7255 8133 7267 8167
rect 7301 8133 7313 8167
rect 7255 8099 7313 8133
rect 7255 8065 7267 8099
rect 7301 8065 7313 8099
rect 7255 8031 7313 8065
rect 7255 7997 7267 8031
rect 7301 7997 7313 8031
rect 7255 7982 7313 7997
rect 7513 8167 7571 8182
rect 7513 8133 7525 8167
rect 7559 8133 7571 8167
rect 7513 8099 7571 8133
rect 7513 8065 7525 8099
rect 7559 8065 7571 8099
rect 7513 8031 7571 8065
rect 7513 7997 7525 8031
rect 7559 7997 7571 8031
rect 7513 7982 7571 7997
rect 7771 8167 7829 8182
rect 7771 8133 7783 8167
rect 7817 8133 7829 8167
rect 7771 8099 7829 8133
rect 7771 8065 7783 8099
rect 7817 8065 7829 8099
rect 7771 8031 7829 8065
rect 7771 7997 7783 8031
rect 7817 7997 7829 8031
rect 7771 7982 7829 7997
rect 8029 8167 8087 8182
rect 8029 8133 8041 8167
rect 8075 8133 8087 8167
rect 8029 8099 8087 8133
rect 8029 8065 8041 8099
rect 8075 8065 8087 8099
rect 8029 8031 8087 8065
rect 8029 7997 8041 8031
rect 8075 7997 8087 8031
rect 8029 7982 8087 7997
rect 8287 8167 8345 8182
rect 8287 8133 8299 8167
rect 8333 8133 8345 8167
rect 8287 8099 8345 8133
rect 8287 8065 8299 8099
rect 8333 8065 8345 8099
rect 8287 8031 8345 8065
rect 8287 7997 8299 8031
rect 8333 7997 8345 8031
rect 8287 7982 8345 7997
rect 8545 8167 8603 8182
rect 8545 8133 8557 8167
rect 8591 8133 8603 8167
rect 8545 8099 8603 8133
rect 8545 8065 8557 8099
rect 8591 8065 8603 8099
rect 8545 8031 8603 8065
rect 8545 7997 8557 8031
rect 8591 7997 8603 8031
rect 8545 7982 8603 7997
<< ndiffc >>
rect 3083 10650 3117 10684
rect 3083 10582 3117 10616
rect 3083 10514 3117 10548
rect 3341 10650 3375 10684
rect 3341 10582 3375 10616
rect 3341 10514 3375 10548
rect 3599 10650 3633 10684
rect 3599 10582 3633 10616
rect 3599 10514 3633 10548
rect 3857 10650 3891 10684
rect 3857 10582 3891 10616
rect 3857 10514 3891 10548
rect 4115 10650 4149 10684
rect 4115 10582 4149 10616
rect 4115 10514 4149 10548
rect 4373 10650 4407 10684
rect 4373 10582 4407 10616
rect 4373 10514 4407 10548
rect 4631 10650 4665 10684
rect 4631 10582 4665 10616
rect 4631 10514 4665 10548
rect 4889 10650 4923 10684
rect 4889 10582 4923 10616
rect 4889 10514 4923 10548
rect 5147 10650 5181 10684
rect 5147 10582 5181 10616
rect 5147 10514 5181 10548
rect 3083 10232 3117 10266
rect 3083 10164 3117 10198
rect 3083 10096 3117 10130
rect 3341 10232 3375 10266
rect 3341 10164 3375 10198
rect 3341 10096 3375 10130
rect 3599 10232 3633 10266
rect 3599 10164 3633 10198
rect 3599 10096 3633 10130
rect 3857 10232 3891 10266
rect 3857 10164 3891 10198
rect 3857 10096 3891 10130
rect 4115 10232 4149 10266
rect 4115 10164 4149 10198
rect 4115 10096 4149 10130
rect 4373 10232 4407 10266
rect 4373 10164 4407 10198
rect 4373 10096 4407 10130
rect 4631 10232 4665 10266
rect 4631 10164 4665 10198
rect 4631 10096 4665 10130
rect 4889 10232 4923 10266
rect 4889 10164 4923 10198
rect 4889 10096 4923 10130
rect 5147 10232 5181 10266
rect 5147 10164 5181 10198
rect 5147 10096 5181 10130
rect 3083 9814 3117 9848
rect 3083 9746 3117 9780
rect 3083 9678 3117 9712
rect 3341 9814 3375 9848
rect 3341 9746 3375 9780
rect 3341 9678 3375 9712
rect 3599 9814 3633 9848
rect 3599 9746 3633 9780
rect 3599 9678 3633 9712
rect 3857 9814 3891 9848
rect 3857 9746 3891 9780
rect 3857 9678 3891 9712
rect 4115 9814 4149 9848
rect 4115 9746 4149 9780
rect 4115 9678 4149 9712
rect 4373 9814 4407 9848
rect 4373 9746 4407 9780
rect 4373 9678 4407 9712
rect 4631 9814 4665 9848
rect 4631 9746 4665 9780
rect 4631 9678 4665 9712
rect 4889 9814 4923 9848
rect 4889 9746 4923 9780
rect 4889 9678 4923 9712
rect 5147 9814 5181 9848
rect 5147 9746 5181 9780
rect 5147 9678 5181 9712
rect 3083 9396 3117 9430
rect 3083 9328 3117 9362
rect 3083 9260 3117 9294
rect 3341 9396 3375 9430
rect 3341 9328 3375 9362
rect 3341 9260 3375 9294
rect 3599 9396 3633 9430
rect 3599 9328 3633 9362
rect 3599 9260 3633 9294
rect 3857 9396 3891 9430
rect 3857 9328 3891 9362
rect 3857 9260 3891 9294
rect 4115 9396 4149 9430
rect 4115 9328 4149 9362
rect 4115 9260 4149 9294
rect 4373 9396 4407 9430
rect 4373 9328 4407 9362
rect 4373 9260 4407 9294
rect 4631 9396 4665 9430
rect 4631 9328 4665 9362
rect 4631 9260 4665 9294
rect 4889 9396 4923 9430
rect 4889 9328 4923 9362
rect 4889 9260 4923 9294
rect 5147 9396 5181 9430
rect 5147 9328 5181 9362
rect 5147 9260 5181 9294
rect 3083 8974 3117 9008
rect 3083 8906 3117 8940
rect 3083 8838 3117 8872
rect 3341 8974 3375 9008
rect 3341 8906 3375 8940
rect 3341 8838 3375 8872
rect 3599 8974 3633 9008
rect 3599 8906 3633 8940
rect 3599 8838 3633 8872
rect 3857 8974 3891 9008
rect 3857 8906 3891 8940
rect 3857 8838 3891 8872
rect 4115 8974 4149 9008
rect 4115 8906 4149 8940
rect 4115 8838 4149 8872
rect 4373 8974 4407 9008
rect 4373 8906 4407 8940
rect 4373 8838 4407 8872
rect 4631 8974 4665 9008
rect 4631 8906 4665 8940
rect 4631 8838 4665 8872
rect 4889 8974 4923 9008
rect 4889 8906 4923 8940
rect 4889 8838 4923 8872
rect 5147 8974 5181 9008
rect 5147 8906 5181 8940
rect 5147 8838 5181 8872
rect 3083 8552 3117 8586
rect 3083 8484 3117 8518
rect 3083 8416 3117 8450
rect 3341 8552 3375 8586
rect 3341 8484 3375 8518
rect 3341 8416 3375 8450
rect 3599 8552 3633 8586
rect 3599 8484 3633 8518
rect 3599 8416 3633 8450
rect 3857 8552 3891 8586
rect 3857 8484 3891 8518
rect 3857 8416 3891 8450
rect 4115 8552 4149 8586
rect 4115 8484 4149 8518
rect 4115 8416 4149 8450
rect 4373 8552 4407 8586
rect 4373 8484 4407 8518
rect 4373 8416 4407 8450
rect 4631 8552 4665 8586
rect 4631 8484 4665 8518
rect 4631 8416 4665 8450
rect 4889 8552 4923 8586
rect 4889 8484 4923 8518
rect 4889 8416 4923 8450
rect 5147 8552 5181 8586
rect 5147 8484 5181 8518
rect 5147 8416 5181 8450
rect -2208 7901 -2174 7935
rect -2208 7833 -2174 7867
rect -2208 7765 -2174 7799
rect -1950 7901 -1916 7935
rect -1950 7833 -1916 7867
rect -1950 7765 -1916 7799
rect -1692 7901 -1658 7935
rect -1692 7833 -1658 7867
rect -1692 7765 -1658 7799
rect -1434 7901 -1400 7935
rect -1434 7833 -1400 7867
rect -1434 7765 -1400 7799
rect -1176 7901 -1142 7935
rect -1176 7833 -1142 7867
rect -1176 7765 -1142 7799
rect -918 7901 -884 7935
rect -918 7833 -884 7867
rect -918 7765 -884 7799
rect -660 7901 -626 7935
rect -660 7833 -626 7867
rect -660 7765 -626 7799
rect -402 7901 -368 7935
rect -402 7833 -368 7867
rect -402 7765 -368 7799
rect -144 7901 -110 7935
rect -144 7833 -110 7867
rect -144 7765 -110 7799
rect 114 7901 148 7935
rect 114 7833 148 7867
rect 114 7765 148 7799
rect 372 7901 406 7935
rect 372 7833 406 7867
rect 372 7765 406 7799
rect 630 7901 664 7935
rect 630 7833 664 7867
rect 630 7765 664 7799
rect 888 7901 922 7935
rect 888 7833 922 7867
rect 888 7765 922 7799
rect 1146 7901 1180 7935
rect 1146 7833 1180 7867
rect 1146 7765 1180 7799
rect 1404 7901 1438 7935
rect 1404 7833 1438 7867
rect 1404 7765 1438 7799
rect -2208 7483 -2174 7517
rect -2208 7415 -2174 7449
rect -2208 7347 -2174 7381
rect -1950 7483 -1916 7517
rect -1950 7415 -1916 7449
rect -1950 7347 -1916 7381
rect -1692 7483 -1658 7517
rect -1692 7415 -1658 7449
rect -1692 7347 -1658 7381
rect -1434 7483 -1400 7517
rect -1434 7415 -1400 7449
rect -1434 7347 -1400 7381
rect -1176 7483 -1142 7517
rect -1176 7415 -1142 7449
rect -1176 7347 -1142 7381
rect -918 7483 -884 7517
rect -918 7415 -884 7449
rect -918 7347 -884 7381
rect -660 7483 -626 7517
rect -660 7415 -626 7449
rect -660 7347 -626 7381
rect -402 7483 -368 7517
rect -402 7415 -368 7449
rect -402 7347 -368 7381
rect -144 7483 -110 7517
rect -144 7415 -110 7449
rect -144 7347 -110 7381
rect 114 7483 148 7517
rect 114 7415 148 7449
rect 114 7347 148 7381
rect 372 7483 406 7517
rect 372 7415 406 7449
rect 372 7347 406 7381
rect 630 7483 664 7517
rect 630 7415 664 7449
rect 630 7347 664 7381
rect 888 7483 922 7517
rect 888 7415 922 7449
rect 888 7347 922 7381
rect 1146 7483 1180 7517
rect 1146 7415 1180 7449
rect 1146 7347 1180 7381
rect 1404 7483 1438 7517
rect 1404 7415 1438 7449
rect 1404 7347 1438 7381
rect -2208 7065 -2174 7099
rect -2208 6997 -2174 7031
rect -2208 6929 -2174 6963
rect -1950 7065 -1916 7099
rect -1950 6997 -1916 7031
rect -1950 6929 -1916 6963
rect -1692 7065 -1658 7099
rect -1692 6997 -1658 7031
rect -1692 6929 -1658 6963
rect -1434 7065 -1400 7099
rect -1434 6997 -1400 7031
rect -1434 6929 -1400 6963
rect -1176 7065 -1142 7099
rect -1176 6997 -1142 7031
rect -1176 6929 -1142 6963
rect -918 7065 -884 7099
rect -918 6997 -884 7031
rect -918 6929 -884 6963
rect -660 7065 -626 7099
rect -660 6997 -626 7031
rect -660 6929 -626 6963
rect -402 7065 -368 7099
rect -402 6997 -368 7031
rect -402 6929 -368 6963
rect -144 7065 -110 7099
rect -144 6997 -110 7031
rect -144 6929 -110 6963
rect 114 7065 148 7099
rect 114 6997 148 7031
rect 114 6929 148 6963
rect 372 7065 406 7099
rect 372 6997 406 7031
rect 372 6929 406 6963
rect 630 7065 664 7099
rect 630 6997 664 7031
rect 630 6929 664 6963
rect 888 7065 922 7099
rect 888 6997 922 7031
rect 888 6929 922 6963
rect 1146 7065 1180 7099
rect 1146 6997 1180 7031
rect 1146 6929 1180 6963
rect 1404 7065 1438 7099
rect 1404 6997 1438 7031
rect 1404 6929 1438 6963
rect -2208 6647 -2174 6681
rect -2208 6579 -2174 6613
rect -2208 6511 -2174 6545
rect -1950 6647 -1916 6681
rect -1950 6579 -1916 6613
rect -1950 6511 -1916 6545
rect -1692 6647 -1658 6681
rect -1692 6579 -1658 6613
rect -1692 6511 -1658 6545
rect -1434 6647 -1400 6681
rect -1434 6579 -1400 6613
rect -1434 6511 -1400 6545
rect -1176 6647 -1142 6681
rect -1176 6579 -1142 6613
rect -1176 6511 -1142 6545
rect -918 6647 -884 6681
rect -918 6579 -884 6613
rect -918 6511 -884 6545
rect -660 6647 -626 6681
rect -660 6579 -626 6613
rect -660 6511 -626 6545
rect -402 6647 -368 6681
rect -402 6579 -368 6613
rect -402 6511 -368 6545
rect -144 6647 -110 6681
rect -144 6579 -110 6613
rect -144 6511 -110 6545
rect 114 6647 148 6681
rect 114 6579 148 6613
rect 114 6511 148 6545
rect 372 6647 406 6681
rect 372 6579 406 6613
rect 372 6511 406 6545
rect 630 6647 664 6681
rect 630 6579 664 6613
rect 630 6511 664 6545
rect 888 6647 922 6681
rect 888 6579 922 6613
rect 888 6511 922 6545
rect 1146 6647 1180 6681
rect 1146 6579 1180 6613
rect 1146 6511 1180 6545
rect 1404 6647 1438 6681
rect 1404 6579 1438 6613
rect 1404 6511 1438 6545
rect -2208 6229 -2174 6263
rect -2208 6161 -2174 6195
rect -2208 6093 -2174 6127
rect -1950 6229 -1916 6263
rect -1950 6161 -1916 6195
rect -1950 6093 -1916 6127
rect -1692 6229 -1658 6263
rect -1692 6161 -1658 6195
rect -1692 6093 -1658 6127
rect -1434 6229 -1400 6263
rect -1434 6161 -1400 6195
rect -1434 6093 -1400 6127
rect -1176 6229 -1142 6263
rect -1176 6161 -1142 6195
rect -1176 6093 -1142 6127
rect -918 6229 -884 6263
rect -918 6161 -884 6195
rect -918 6093 -884 6127
rect -660 6229 -626 6263
rect -660 6161 -626 6195
rect -660 6093 -626 6127
rect -402 6229 -368 6263
rect -402 6161 -368 6195
rect -402 6093 -368 6127
rect -144 6229 -110 6263
rect -144 6161 -110 6195
rect -144 6093 -110 6127
rect 114 6229 148 6263
rect 114 6161 148 6195
rect 114 6093 148 6127
rect 372 6229 406 6263
rect 372 6161 406 6195
rect 372 6093 406 6127
rect 630 6229 664 6263
rect 630 6161 664 6195
rect 630 6093 664 6127
rect 888 6229 922 6263
rect 888 6161 922 6195
rect 888 6093 922 6127
rect 1146 6229 1180 6263
rect 1146 6161 1180 6195
rect 1146 6093 1180 6127
rect 1404 6229 1438 6263
rect 1404 6161 1438 6195
rect 1404 6093 1438 6127
rect -2208 5811 -2174 5845
rect -2208 5743 -2174 5777
rect -2208 5675 -2174 5709
rect -1950 5811 -1916 5845
rect -1950 5743 -1916 5777
rect -1950 5675 -1916 5709
rect -1692 5811 -1658 5845
rect -1692 5743 -1658 5777
rect -1692 5675 -1658 5709
rect -1434 5811 -1400 5845
rect -1434 5743 -1400 5777
rect -1434 5675 -1400 5709
rect -1176 5811 -1142 5845
rect -1176 5743 -1142 5777
rect -1176 5675 -1142 5709
rect -918 5811 -884 5845
rect -918 5743 -884 5777
rect -918 5675 -884 5709
rect -660 5811 -626 5845
rect -660 5743 -626 5777
rect -660 5675 -626 5709
rect -402 5811 -368 5845
rect -402 5743 -368 5777
rect -402 5675 -368 5709
rect -144 5811 -110 5845
rect -144 5743 -110 5777
rect -144 5675 -110 5709
rect 114 5811 148 5845
rect 114 5743 148 5777
rect 114 5675 148 5709
rect 372 5811 406 5845
rect 372 5743 406 5777
rect 372 5675 406 5709
rect 630 5811 664 5845
rect 630 5743 664 5777
rect 630 5675 664 5709
rect 888 5811 922 5845
rect 888 5743 922 5777
rect 888 5675 922 5709
rect 1146 5811 1180 5845
rect 1146 5743 1180 5777
rect 1146 5675 1180 5709
rect 1404 5811 1438 5845
rect 1404 5743 1438 5777
rect 1404 5675 1438 5709
rect -2208 5393 -2174 5427
rect -2208 5325 -2174 5359
rect -2208 5257 -2174 5291
rect -1950 5393 -1916 5427
rect -1950 5325 -1916 5359
rect -1950 5257 -1916 5291
rect -1692 5393 -1658 5427
rect -1692 5325 -1658 5359
rect -1692 5257 -1658 5291
rect -1434 5393 -1400 5427
rect -1434 5325 -1400 5359
rect -1434 5257 -1400 5291
rect -1176 5393 -1142 5427
rect -1176 5325 -1142 5359
rect -1176 5257 -1142 5291
rect -918 5393 -884 5427
rect -918 5325 -884 5359
rect -918 5257 -884 5291
rect -660 5393 -626 5427
rect -660 5325 -626 5359
rect -660 5257 -626 5291
rect -402 5393 -368 5427
rect -402 5325 -368 5359
rect -402 5257 -368 5291
rect -144 5393 -110 5427
rect -144 5325 -110 5359
rect -144 5257 -110 5291
rect 114 5393 148 5427
rect 114 5325 148 5359
rect 114 5257 148 5291
rect 372 5393 406 5427
rect 372 5325 406 5359
rect 372 5257 406 5291
rect 630 5393 664 5427
rect 630 5325 664 5359
rect 630 5257 664 5291
rect 888 5393 922 5427
rect 888 5325 922 5359
rect 888 5257 922 5291
rect 1146 5393 1180 5427
rect 1146 5325 1180 5359
rect 1146 5257 1180 5291
rect 1404 5393 1438 5427
rect 1404 5325 1438 5359
rect 1404 5257 1438 5291
rect -2208 4975 -2174 5009
rect -2208 4907 -2174 4941
rect -2208 4839 -2174 4873
rect -1950 4975 -1916 5009
rect -1950 4907 -1916 4941
rect -1950 4839 -1916 4873
rect -1692 4975 -1658 5009
rect -1692 4907 -1658 4941
rect -1692 4839 -1658 4873
rect -1434 4975 -1400 5009
rect -1434 4907 -1400 4941
rect -1434 4839 -1400 4873
rect -1176 4975 -1142 5009
rect -1176 4907 -1142 4941
rect -1176 4839 -1142 4873
rect -918 4975 -884 5009
rect -918 4907 -884 4941
rect -918 4839 -884 4873
rect -660 4975 -626 5009
rect -660 4907 -626 4941
rect -660 4839 -626 4873
rect -402 4975 -368 5009
rect -402 4907 -368 4941
rect -402 4839 -368 4873
rect -144 4975 -110 5009
rect -144 4907 -110 4941
rect -144 4839 -110 4873
rect 114 4975 148 5009
rect 114 4907 148 4941
rect 114 4839 148 4873
rect 372 4975 406 5009
rect 372 4907 406 4941
rect 372 4839 406 4873
rect 630 4975 664 5009
rect 630 4907 664 4941
rect 630 4839 664 4873
rect 888 4975 922 5009
rect 888 4907 922 4941
rect 888 4839 922 4873
rect 1146 4975 1180 5009
rect 1146 4907 1180 4941
rect 1146 4839 1180 4873
rect 1404 4975 1438 5009
rect 1404 4907 1438 4941
rect 1404 4839 1438 4873
rect -2208 4557 -2174 4591
rect -2208 4489 -2174 4523
rect -2208 4421 -2174 4455
rect -1950 4557 -1916 4591
rect -1950 4489 -1916 4523
rect -1950 4421 -1916 4455
rect -1692 4557 -1658 4591
rect -1692 4489 -1658 4523
rect -1692 4421 -1658 4455
rect -1434 4557 -1400 4591
rect -1434 4489 -1400 4523
rect -1434 4421 -1400 4455
rect -1176 4557 -1142 4591
rect -1176 4489 -1142 4523
rect -1176 4421 -1142 4455
rect -918 4557 -884 4591
rect -918 4489 -884 4523
rect -918 4421 -884 4455
rect -660 4557 -626 4591
rect -660 4489 -626 4523
rect -660 4421 -626 4455
rect -402 4557 -368 4591
rect -402 4489 -368 4523
rect -402 4421 -368 4455
rect -144 4557 -110 4591
rect -144 4489 -110 4523
rect -144 4421 -110 4455
rect 114 4557 148 4591
rect 114 4489 148 4523
rect 114 4421 148 4455
rect 372 4557 406 4591
rect 372 4489 406 4523
rect 372 4421 406 4455
rect 630 4557 664 4591
rect 630 4489 664 4523
rect 630 4421 664 4455
rect 888 4557 922 4591
rect 888 4489 922 4523
rect 888 4421 922 4455
rect 1146 4557 1180 4591
rect 1146 4489 1180 4523
rect 1146 4421 1180 4455
rect 1404 4557 1438 4591
rect 1404 4489 1438 4523
rect 1404 4421 1438 4455
rect -2208 4139 -2174 4173
rect -2208 4071 -2174 4105
rect -2208 4003 -2174 4037
rect -1950 4139 -1916 4173
rect -1950 4071 -1916 4105
rect -1950 4003 -1916 4037
rect -1692 4139 -1658 4173
rect -1692 4071 -1658 4105
rect -1692 4003 -1658 4037
rect -1434 4139 -1400 4173
rect -1434 4071 -1400 4105
rect -1434 4003 -1400 4037
rect -1176 4139 -1142 4173
rect -1176 4071 -1142 4105
rect -1176 4003 -1142 4037
rect -918 4139 -884 4173
rect -918 4071 -884 4105
rect -918 4003 -884 4037
rect -660 4139 -626 4173
rect -660 4071 -626 4105
rect -660 4003 -626 4037
rect -402 4139 -368 4173
rect -402 4071 -368 4105
rect -402 4003 -368 4037
rect -144 4139 -110 4173
rect -144 4071 -110 4105
rect -144 4003 -110 4037
rect 114 4139 148 4173
rect 114 4071 148 4105
rect 114 4003 148 4037
rect 372 4139 406 4173
rect 372 4071 406 4105
rect 372 4003 406 4037
rect 630 4139 664 4173
rect 630 4071 664 4105
rect 630 4003 664 4037
rect 888 4139 922 4173
rect 888 4071 922 4105
rect 888 4003 922 4037
rect 1146 4139 1180 4173
rect 1146 4071 1180 4105
rect 1146 4003 1180 4037
rect 1404 4139 1438 4173
rect 1404 4071 1438 4105
rect 1404 4003 1438 4037
rect 3622 7262 3656 7296
rect 3622 7194 3656 7228
rect 3622 7126 3656 7160
rect 3880 7262 3914 7296
rect 3880 7194 3914 7228
rect 3880 7126 3914 7160
rect 4138 7262 4172 7296
rect 4138 7194 4172 7228
rect 4138 7126 4172 7160
rect 4396 7262 4430 7296
rect 4396 7194 4430 7228
rect 4396 7126 4430 7160
rect 4654 7262 4688 7296
rect 4654 7194 4688 7228
rect 4654 7126 4688 7160
rect 4912 7262 4946 7296
rect 4912 7194 4946 7228
rect 4912 7126 4946 7160
rect 5170 7262 5204 7296
rect 5170 7194 5204 7228
rect 5170 7126 5204 7160
rect 5428 7262 5462 7296
rect 5428 7194 5462 7228
rect 5428 7126 5462 7160
rect 5686 7262 5720 7296
rect 5686 7194 5720 7228
rect 5686 7126 5720 7160
rect 5944 7262 5978 7296
rect 5944 7194 5978 7228
rect 5944 7126 5978 7160
rect 6202 7262 6236 7296
rect 6202 7194 6236 7228
rect 6202 7126 6236 7160
rect 3622 6844 3656 6878
rect 3622 6776 3656 6810
rect 3622 6708 3656 6742
rect 3880 6844 3914 6878
rect 3880 6776 3914 6810
rect 3880 6708 3914 6742
rect 4138 6844 4172 6878
rect 4138 6776 4172 6810
rect 4138 6708 4172 6742
rect 4396 6844 4430 6878
rect 4396 6776 4430 6810
rect 4396 6708 4430 6742
rect 4654 6844 4688 6878
rect 4654 6776 4688 6810
rect 4654 6708 4688 6742
rect 4912 6844 4946 6878
rect 4912 6776 4946 6810
rect 4912 6708 4946 6742
rect 5170 6844 5204 6878
rect 5170 6776 5204 6810
rect 5170 6708 5204 6742
rect 5428 6844 5462 6878
rect 5428 6776 5462 6810
rect 5428 6708 5462 6742
rect 5686 6844 5720 6878
rect 5686 6776 5720 6810
rect 5686 6708 5720 6742
rect 5944 6844 5978 6878
rect 5944 6776 5978 6810
rect 5944 6708 5978 6742
rect 6202 6844 6236 6878
rect 6202 6776 6236 6810
rect 6202 6708 6236 6742
rect 3622 6426 3656 6460
rect 3622 6358 3656 6392
rect 3622 6290 3656 6324
rect 3880 6426 3914 6460
rect 3880 6358 3914 6392
rect 3880 6290 3914 6324
rect 4138 6426 4172 6460
rect 4138 6358 4172 6392
rect 4138 6290 4172 6324
rect 4396 6426 4430 6460
rect 4396 6358 4430 6392
rect 4396 6290 4430 6324
rect 4654 6426 4688 6460
rect 4654 6358 4688 6392
rect 4654 6290 4688 6324
rect 4912 6426 4946 6460
rect 4912 6358 4946 6392
rect 4912 6290 4946 6324
rect 5170 6426 5204 6460
rect 5170 6358 5204 6392
rect 5170 6290 5204 6324
rect 5428 6426 5462 6460
rect 5428 6358 5462 6392
rect 5428 6290 5462 6324
rect 5686 6426 5720 6460
rect 5686 6358 5720 6392
rect 5686 6290 5720 6324
rect 5944 6426 5978 6460
rect 5944 6358 5978 6392
rect 5944 6290 5978 6324
rect 6202 6426 6236 6460
rect 6202 6358 6236 6392
rect 6202 6290 6236 6324
rect 3622 6008 3656 6042
rect 3622 5940 3656 5974
rect 3622 5872 3656 5906
rect 3880 6008 3914 6042
rect 3880 5940 3914 5974
rect 3880 5872 3914 5906
rect 4138 6008 4172 6042
rect 4138 5940 4172 5974
rect 4138 5872 4172 5906
rect 4396 6008 4430 6042
rect 4396 5940 4430 5974
rect 4396 5872 4430 5906
rect 4654 6008 4688 6042
rect 4654 5940 4688 5974
rect 4654 5872 4688 5906
rect 4912 6008 4946 6042
rect 4912 5940 4946 5974
rect 4912 5872 4946 5906
rect 5170 6008 5204 6042
rect 5170 5940 5204 5974
rect 5170 5872 5204 5906
rect 5428 6008 5462 6042
rect 5428 5940 5462 5974
rect 5428 5872 5462 5906
rect 5686 6008 5720 6042
rect 5686 5940 5720 5974
rect 5686 5872 5720 5906
rect 5944 6008 5978 6042
rect 5944 5940 5978 5974
rect 5944 5872 5978 5906
rect 6202 6008 6236 6042
rect 6202 5940 6236 5974
rect 6202 5872 6236 5906
rect 3622 5590 3656 5624
rect 3622 5522 3656 5556
rect 3622 5454 3656 5488
rect 3880 5590 3914 5624
rect 3880 5522 3914 5556
rect 3880 5454 3914 5488
rect 4138 5590 4172 5624
rect 4138 5522 4172 5556
rect 4138 5454 4172 5488
rect 4396 5590 4430 5624
rect 4396 5522 4430 5556
rect 4396 5454 4430 5488
rect 4654 5590 4688 5624
rect 4654 5522 4688 5556
rect 4654 5454 4688 5488
rect 4912 5590 4946 5624
rect 4912 5522 4946 5556
rect 4912 5454 4946 5488
rect 5170 5590 5204 5624
rect 5170 5522 5204 5556
rect 5170 5454 5204 5488
rect 5428 5590 5462 5624
rect 5428 5522 5462 5556
rect 5428 5454 5462 5488
rect 5686 5590 5720 5624
rect 5686 5522 5720 5556
rect 5686 5454 5720 5488
rect 5944 5590 5978 5624
rect 5944 5522 5978 5556
rect 5944 5454 5978 5488
rect 6202 5590 6236 5624
rect 6202 5522 6236 5556
rect 6202 5454 6236 5488
rect 3622 5172 3656 5206
rect 3622 5104 3656 5138
rect 3622 5036 3656 5070
rect 3880 5172 3914 5206
rect 3880 5104 3914 5138
rect 3880 5036 3914 5070
rect 4138 5172 4172 5206
rect 4138 5104 4172 5138
rect 4138 5036 4172 5070
rect 4396 5172 4430 5206
rect 4396 5104 4430 5138
rect 4396 5036 4430 5070
rect 4654 5172 4688 5206
rect 4654 5104 4688 5138
rect 4654 5036 4688 5070
rect 4912 5172 4946 5206
rect 4912 5104 4946 5138
rect 4912 5036 4946 5070
rect 5170 5172 5204 5206
rect 5170 5104 5204 5138
rect 5170 5036 5204 5070
rect 5428 5172 5462 5206
rect 5428 5104 5462 5138
rect 5428 5036 5462 5070
rect 5686 5172 5720 5206
rect 5686 5104 5720 5138
rect 5686 5036 5720 5070
rect 5944 5172 5978 5206
rect 5944 5104 5978 5138
rect 5944 5036 5978 5070
rect 6202 5172 6236 5206
rect 6202 5104 6236 5138
rect 6202 5036 6236 5070
rect 3622 4754 3656 4788
rect 3622 4686 3656 4720
rect 3622 4618 3656 4652
rect 3880 4754 3914 4788
rect 3880 4686 3914 4720
rect 3880 4618 3914 4652
rect 4138 4754 4172 4788
rect 4138 4686 4172 4720
rect 4138 4618 4172 4652
rect 4396 4754 4430 4788
rect 4396 4686 4430 4720
rect 4396 4618 4430 4652
rect 4654 4754 4688 4788
rect 4654 4686 4688 4720
rect 4654 4618 4688 4652
rect 4912 4754 4946 4788
rect 4912 4686 4946 4720
rect 4912 4618 4946 4652
rect 5170 4754 5204 4788
rect 5170 4686 5204 4720
rect 5170 4618 5204 4652
rect 5428 4754 5462 4788
rect 5428 4686 5462 4720
rect 5428 4618 5462 4652
rect 5686 4754 5720 4788
rect 5686 4686 5720 4720
rect 5686 4618 5720 4652
rect 5944 4754 5978 4788
rect 5944 4686 5978 4720
rect 5944 4618 5978 4652
rect 6202 4754 6236 4788
rect 6202 4686 6236 4720
rect 6202 4618 6236 4652
rect 3622 4336 3656 4370
rect 3622 4268 3656 4302
rect 3622 4200 3656 4234
rect 3880 4336 3914 4370
rect 3880 4268 3914 4302
rect 3880 4200 3914 4234
rect 4138 4336 4172 4370
rect 4138 4268 4172 4302
rect 4138 4200 4172 4234
rect 4396 4336 4430 4370
rect 4396 4268 4430 4302
rect 4396 4200 4430 4234
rect 4654 4336 4688 4370
rect 4654 4268 4688 4302
rect 4654 4200 4688 4234
rect 4912 4336 4946 4370
rect 4912 4268 4946 4302
rect 4912 4200 4946 4234
rect 5170 4336 5204 4370
rect 5170 4268 5204 4302
rect 5170 4200 5204 4234
rect 5428 4336 5462 4370
rect 5428 4268 5462 4302
rect 5428 4200 5462 4234
rect 5686 4336 5720 4370
rect 5686 4268 5720 4302
rect 5686 4200 5720 4234
rect 5944 4336 5978 4370
rect 5944 4268 5978 4302
rect 5944 4200 5978 4234
rect 6202 4336 6236 4370
rect 6202 4268 6236 4302
rect 6202 4200 6236 4234
rect 8358 6851 8392 6885
rect 8358 6783 8392 6817
rect 8358 6715 8392 6749
rect 8616 6851 8650 6885
rect 8616 6783 8650 6817
rect 8616 6715 8650 6749
rect 8874 6851 8908 6885
rect 8874 6783 8908 6817
rect 8874 6715 8908 6749
rect 9132 6851 9166 6885
rect 9132 6783 9166 6817
rect 9132 6715 9166 6749
rect 9390 6851 9424 6885
rect 9390 6783 9424 6817
rect 9390 6715 9424 6749
rect 9648 6851 9682 6885
rect 9648 6783 9682 6817
rect 9648 6715 9682 6749
rect 9906 6851 9940 6885
rect 9906 6783 9940 6817
rect 9906 6715 9940 6749
rect 8358 6433 8392 6467
rect 8358 6365 8392 6399
rect 8358 6297 8392 6331
rect 8616 6433 8650 6467
rect 8616 6365 8650 6399
rect 8616 6297 8650 6331
rect 8874 6433 8908 6467
rect 8874 6365 8908 6399
rect 8874 6297 8908 6331
rect 9132 6433 9166 6467
rect 9132 6365 9166 6399
rect 9132 6297 9166 6331
rect 9390 6433 9424 6467
rect 9390 6365 9424 6399
rect 9390 6297 9424 6331
rect 9648 6433 9682 6467
rect 9648 6365 9682 6399
rect 9648 6297 9682 6331
rect 9906 6433 9940 6467
rect 9906 6365 9940 6399
rect 9906 6297 9940 6331
rect 8358 6015 8392 6049
rect 8358 5947 8392 5981
rect 8358 5879 8392 5913
rect 8616 6015 8650 6049
rect 8616 5947 8650 5981
rect 8616 5879 8650 5913
rect 8874 6015 8908 6049
rect 8874 5947 8908 5981
rect 8874 5879 8908 5913
rect 9132 6015 9166 6049
rect 9132 5947 9166 5981
rect 9132 5879 9166 5913
rect 9390 6015 9424 6049
rect 9390 5947 9424 5981
rect 9390 5879 9424 5913
rect 9648 6015 9682 6049
rect 9648 5947 9682 5981
rect 9648 5879 9682 5913
rect 9906 6015 9940 6049
rect 9906 5947 9940 5981
rect 9906 5879 9940 5913
rect 8358 5597 8392 5631
rect 8358 5529 8392 5563
rect 8358 5461 8392 5495
rect 8616 5597 8650 5631
rect 8616 5529 8650 5563
rect 8616 5461 8650 5495
rect 8874 5597 8908 5631
rect 8874 5529 8908 5563
rect 8874 5461 8908 5495
rect 9132 5597 9166 5631
rect 9132 5529 9166 5563
rect 9132 5461 9166 5495
rect 9390 5597 9424 5631
rect 9390 5529 9424 5563
rect 9390 5461 9424 5495
rect 9648 5597 9682 5631
rect 9648 5529 9682 5563
rect 9648 5461 9682 5495
rect 9906 5597 9940 5631
rect 9906 5529 9940 5563
rect 9906 5461 9940 5495
rect 8358 5179 8392 5213
rect 8358 5111 8392 5145
rect 8358 5043 8392 5077
rect 8616 5179 8650 5213
rect 8616 5111 8650 5145
rect 8616 5043 8650 5077
rect 8874 5179 8908 5213
rect 8874 5111 8908 5145
rect 8874 5043 8908 5077
rect 9132 5179 9166 5213
rect 9132 5111 9166 5145
rect 9132 5043 9166 5077
rect 9390 5179 9424 5213
rect 9390 5111 9424 5145
rect 9390 5043 9424 5077
rect 9648 5179 9682 5213
rect 9648 5111 9682 5145
rect 9648 5043 9682 5077
rect 9906 5179 9940 5213
rect 9906 5111 9940 5145
rect 9906 5043 9940 5077
rect 8358 4761 8392 4795
rect 8358 4693 8392 4727
rect 8358 4625 8392 4659
rect 8616 4761 8650 4795
rect 8616 4693 8650 4727
rect 8616 4625 8650 4659
rect 8874 4761 8908 4795
rect 8874 4693 8908 4727
rect 8874 4625 8908 4659
rect 9132 4761 9166 4795
rect 9132 4693 9166 4727
rect 9132 4625 9166 4659
rect 9390 4761 9424 4795
rect 9390 4693 9424 4727
rect 9390 4625 9424 4659
rect 9648 4761 9682 4795
rect 9648 4693 9682 4727
rect 9648 4625 9682 4659
rect 9906 4761 9940 4795
rect 9906 4693 9940 4727
rect 9906 4625 9940 4659
rect 8358 4343 8392 4377
rect 8358 4275 8392 4309
rect 8358 4207 8392 4241
rect 8616 4343 8650 4377
rect 8616 4275 8650 4309
rect 8616 4207 8650 4241
rect 8874 4343 8908 4377
rect 8874 4275 8908 4309
rect 8874 4207 8908 4241
rect 9132 4343 9166 4377
rect 9132 4275 9166 4309
rect 9132 4207 9166 4241
rect 9390 4343 9424 4377
rect 9390 4275 9424 4309
rect 9390 4207 9424 4241
rect 9648 4343 9682 4377
rect 9648 4275 9682 4309
rect 9648 4207 9682 4241
rect 9906 4343 9940 4377
rect 9906 4275 9940 4309
rect 9906 4207 9940 4241
<< pdiffc >>
rect -1239 10431 -1205 10465
rect -1239 10363 -1205 10397
rect -1239 10295 -1205 10329
rect -981 10431 -947 10465
rect -981 10363 -947 10397
rect -981 10295 -947 10329
rect -723 10431 -689 10465
rect -723 10363 -689 10397
rect -723 10295 -689 10329
rect -465 10431 -431 10465
rect -465 10363 -431 10397
rect -465 10295 -431 10329
rect -207 10431 -173 10465
rect -207 10363 -173 10397
rect -207 10295 -173 10329
rect 51 10431 85 10465
rect 51 10363 85 10397
rect 51 10295 85 10329
rect 309 10431 343 10465
rect 309 10363 343 10397
rect 309 10295 343 10329
rect -1239 9995 -1205 10029
rect -1239 9927 -1205 9961
rect -1239 9859 -1205 9893
rect -981 9995 -947 10029
rect -981 9927 -947 9961
rect -981 9859 -947 9893
rect -723 9995 -689 10029
rect -723 9927 -689 9961
rect -723 9859 -689 9893
rect -465 9995 -431 10029
rect -465 9927 -431 9961
rect -465 9859 -431 9893
rect -207 9995 -173 10029
rect -207 9927 -173 9961
rect -207 9859 -173 9893
rect 51 9995 85 10029
rect 51 9927 85 9961
rect 51 9859 85 9893
rect 309 9995 343 10029
rect 309 9927 343 9961
rect 309 9859 343 9893
rect -1239 9559 -1205 9593
rect -1239 9491 -1205 9525
rect -1239 9423 -1205 9457
rect -981 9559 -947 9593
rect -981 9491 -947 9525
rect -981 9423 -947 9457
rect -723 9559 -689 9593
rect -723 9491 -689 9525
rect -723 9423 -689 9457
rect -465 9559 -431 9593
rect -465 9491 -431 9525
rect -465 9423 -431 9457
rect -207 9559 -173 9593
rect -207 9491 -173 9525
rect -207 9423 -173 9457
rect 51 9559 85 9593
rect 51 9491 85 9525
rect 51 9423 85 9457
rect 309 9559 343 9593
rect 309 9491 343 9525
rect 309 9423 343 9457
rect -1239 9123 -1205 9157
rect -1239 9055 -1205 9089
rect -1239 8987 -1205 9021
rect -981 9123 -947 9157
rect -981 9055 -947 9089
rect -981 8987 -947 9021
rect -723 9123 -689 9157
rect -723 9055 -689 9089
rect -723 8987 -689 9021
rect -465 9123 -431 9157
rect -465 9055 -431 9089
rect -465 8987 -431 9021
rect -207 9123 -173 9157
rect -207 9055 -173 9089
rect -207 8987 -173 9021
rect 51 9123 85 9157
rect 51 9055 85 9089
rect 51 8987 85 9021
rect 309 9123 343 9157
rect 309 9055 343 9089
rect 309 8987 343 9021
rect 7009 10749 7043 10783
rect 7009 10681 7043 10715
rect 7009 10613 7043 10647
rect 7267 10749 7301 10783
rect 7267 10681 7301 10715
rect 7267 10613 7301 10647
rect 7525 10749 7559 10783
rect 7525 10681 7559 10715
rect 7525 10613 7559 10647
rect 7783 10749 7817 10783
rect 7783 10681 7817 10715
rect 7783 10613 7817 10647
rect 8041 10749 8075 10783
rect 8041 10681 8075 10715
rect 8041 10613 8075 10647
rect 8299 10749 8333 10783
rect 8299 10681 8333 10715
rect 8299 10613 8333 10647
rect 8557 10749 8591 10783
rect 8557 10681 8591 10715
rect 8557 10613 8591 10647
rect 7009 10313 7043 10347
rect 7009 10245 7043 10279
rect 7009 10177 7043 10211
rect 7267 10313 7301 10347
rect 7267 10245 7301 10279
rect 7267 10177 7301 10211
rect 7525 10313 7559 10347
rect 7525 10245 7559 10279
rect 7525 10177 7559 10211
rect 7783 10313 7817 10347
rect 7783 10245 7817 10279
rect 7783 10177 7817 10211
rect 8041 10313 8075 10347
rect 8041 10245 8075 10279
rect 8041 10177 8075 10211
rect 8299 10313 8333 10347
rect 8299 10245 8333 10279
rect 8299 10177 8333 10211
rect 8557 10313 8591 10347
rect 8557 10245 8591 10279
rect 8557 10177 8591 10211
rect 7009 9877 7043 9911
rect 7009 9809 7043 9843
rect 7009 9741 7043 9775
rect 7267 9877 7301 9911
rect 7267 9809 7301 9843
rect 7267 9741 7301 9775
rect 7525 9877 7559 9911
rect 7525 9809 7559 9843
rect 7525 9741 7559 9775
rect 7783 9877 7817 9911
rect 7783 9809 7817 9843
rect 7783 9741 7817 9775
rect 8041 9877 8075 9911
rect 8041 9809 8075 9843
rect 8041 9741 8075 9775
rect 8299 9877 8333 9911
rect 8299 9809 8333 9843
rect 8299 9741 8333 9775
rect 8557 9877 8591 9911
rect 8557 9809 8591 9843
rect 8557 9741 8591 9775
rect 7009 9441 7043 9475
rect 7009 9373 7043 9407
rect 7009 9305 7043 9339
rect 7267 9441 7301 9475
rect 7267 9373 7301 9407
rect 7267 9305 7301 9339
rect 7525 9441 7559 9475
rect 7525 9373 7559 9407
rect 7525 9305 7559 9339
rect 7783 9441 7817 9475
rect 7783 9373 7817 9407
rect 7783 9305 7817 9339
rect 8041 9441 8075 9475
rect 8041 9373 8075 9407
rect 8041 9305 8075 9339
rect 8299 9441 8333 9475
rect 8299 9373 8333 9407
rect 8299 9305 8333 9339
rect 8557 9441 8591 9475
rect 8557 9373 8591 9407
rect 8557 9305 8591 9339
rect 7009 9005 7043 9039
rect 7009 8937 7043 8971
rect 7009 8869 7043 8903
rect 7267 9005 7301 9039
rect 7267 8937 7301 8971
rect 7267 8869 7301 8903
rect 7525 9005 7559 9039
rect 7525 8937 7559 8971
rect 7525 8869 7559 8903
rect 7783 9005 7817 9039
rect 7783 8937 7817 8971
rect 7783 8869 7817 8903
rect 8041 9005 8075 9039
rect 8041 8937 8075 8971
rect 8041 8869 8075 8903
rect 8299 9005 8333 9039
rect 8299 8937 8333 8971
rect 8299 8869 8333 8903
rect 8557 9005 8591 9039
rect 8557 8937 8591 8971
rect 8557 8869 8591 8903
rect 7009 8569 7043 8603
rect 7009 8501 7043 8535
rect 7009 8433 7043 8467
rect 7267 8569 7301 8603
rect 7267 8501 7301 8535
rect 7267 8433 7301 8467
rect 7525 8569 7559 8603
rect 7525 8501 7559 8535
rect 7525 8433 7559 8467
rect 7783 8569 7817 8603
rect 7783 8501 7817 8535
rect 7783 8433 7817 8467
rect 8041 8569 8075 8603
rect 8041 8501 8075 8535
rect 8041 8433 8075 8467
rect 8299 8569 8333 8603
rect 8299 8501 8333 8535
rect 8299 8433 8333 8467
rect 8557 8569 8591 8603
rect 8557 8501 8591 8535
rect 8557 8433 8591 8467
rect 7009 8133 7043 8167
rect 7009 8065 7043 8099
rect 7009 7997 7043 8031
rect 7267 8133 7301 8167
rect 7267 8065 7301 8099
rect 7267 7997 7301 8031
rect 7525 8133 7559 8167
rect 7525 8065 7559 8099
rect 7525 7997 7559 8031
rect 7783 8133 7817 8167
rect 7783 8065 7817 8099
rect 7783 7997 7817 8031
rect 8041 8133 8075 8167
rect 8041 8065 8075 8099
rect 8041 7997 8075 8031
rect 8299 8133 8333 8167
rect 8299 8065 8333 8099
rect 8299 7997 8333 8031
rect 8557 8133 8591 8167
rect 8557 8065 8591 8099
rect 8557 7997 8591 8031
<< psubdiff >>
rect 2969 10839 3089 10873
rect 3123 10839 3157 10873
rect 3191 10839 3225 10873
rect 3259 10839 3293 10873
rect 3327 10839 3361 10873
rect 3395 10839 3429 10873
rect 3463 10839 3497 10873
rect 3531 10839 3565 10873
rect 3599 10839 3633 10873
rect 3667 10839 3701 10873
rect 3735 10839 3769 10873
rect 3803 10839 3837 10873
rect 3871 10839 3905 10873
rect 3939 10839 3973 10873
rect 4007 10839 4041 10873
rect 4075 10839 4109 10873
rect 4143 10839 4177 10873
rect 4211 10839 4245 10873
rect 4279 10839 4313 10873
rect 4347 10839 4381 10873
rect 4415 10839 4449 10873
rect 4483 10839 4517 10873
rect 4551 10839 4585 10873
rect 4619 10839 4653 10873
rect 4687 10839 4721 10873
rect 4755 10839 4789 10873
rect 4823 10839 4857 10873
rect 4891 10839 4925 10873
rect 4959 10839 4993 10873
rect 5027 10839 5061 10873
rect 5095 10839 5129 10873
rect 5163 10839 5296 10873
rect 2969 10771 3003 10839
rect 2969 10703 3003 10737
rect 5262 10771 5296 10839
rect 5262 10703 5296 10737
rect 2969 10635 3003 10669
rect 2969 10567 3003 10601
rect 2969 10499 3003 10533
rect 5262 10635 5296 10669
rect 5262 10567 5296 10601
rect 5262 10499 5296 10533
rect 2969 10431 3003 10465
rect 5262 10431 5296 10465
rect 2969 10363 3003 10397
rect 2969 10295 3003 10329
rect 5262 10363 5296 10397
rect 5262 10295 5296 10329
rect 2969 10227 3003 10261
rect 2969 10159 3003 10193
rect 2969 10091 3003 10125
rect 5262 10227 5296 10261
rect 5262 10159 5296 10193
rect 5262 10091 5296 10125
rect 2969 10023 3003 10057
rect 5262 10023 5296 10057
rect 2969 9955 3003 9989
rect 5262 9955 5296 9989
rect 2969 9887 3003 9921
rect 5262 9887 5296 9921
rect 2969 9819 3003 9853
rect 2969 9751 3003 9785
rect 2969 9683 3003 9717
rect 5262 9819 5296 9853
rect 5262 9751 5296 9785
rect 5262 9683 5296 9717
rect 2969 9615 3003 9649
rect 2969 9547 3003 9581
rect 5262 9615 5296 9649
rect 5262 9547 5296 9581
rect 2969 9479 3003 9513
rect 5262 9479 5296 9513
rect 2969 9411 3003 9445
rect 2969 9343 3003 9377
rect 2969 9275 3003 9309
rect 5262 9411 5296 9445
rect 5262 9343 5296 9377
rect 5262 9275 5296 9309
rect 2969 9207 3003 9241
rect 2969 9139 3003 9173
rect 5262 9207 5296 9241
rect 5262 9139 5296 9173
rect 2969 9071 3003 9105
rect 2969 9003 3003 9037
rect 5262 9071 5296 9105
rect 2969 8935 3003 8969
rect 2969 8867 3003 8901
rect 2969 8799 3003 8833
rect 5262 9003 5296 9037
rect 5262 8935 5296 8969
rect 5262 8867 5296 8901
rect 2969 8731 3003 8765
rect 5262 8799 5296 8833
rect 2969 8663 3003 8697
rect 5262 8731 5296 8765
rect 2969 8595 3003 8629
rect 5262 8663 5296 8697
rect 2969 8527 3003 8561
rect 2969 8459 3003 8493
rect 2969 8391 3003 8425
rect 5262 8595 5296 8629
rect 5262 8527 5296 8561
rect 5262 8459 5296 8493
rect 2969 8268 3003 8357
rect 5262 8391 5296 8425
rect 5262 8268 5296 8357
rect 2969 8234 3089 8268
rect 3123 8234 3157 8268
rect 3191 8234 3225 8268
rect 3259 8234 3293 8268
rect 3327 8234 3361 8268
rect 3395 8234 3429 8268
rect 3463 8234 3497 8268
rect 3531 8234 3565 8268
rect 3599 8234 3633 8268
rect 3667 8234 3701 8268
rect 3735 8234 3769 8268
rect 3803 8234 3837 8268
rect 3871 8234 3905 8268
rect 3939 8234 3973 8268
rect 4007 8234 4041 8268
rect 4075 8234 4109 8268
rect 4143 8234 4177 8268
rect 4211 8234 4245 8268
rect 4279 8234 4313 8268
rect 4347 8234 4381 8268
rect 4415 8234 4449 8268
rect 4483 8234 4517 8268
rect 4551 8234 4585 8268
rect 4619 8234 4653 8268
rect 4687 8234 4721 8268
rect 4755 8234 4789 8268
rect 4823 8234 4857 8268
rect 4891 8234 4925 8268
rect 4959 8234 4993 8268
rect 5027 8234 5061 8268
rect 5095 8234 5129 8268
rect 5163 8234 5296 8268
rect -2322 8090 -2202 8124
rect -2168 8090 -2134 8124
rect -2100 8090 -2066 8124
rect -2032 8090 -1998 8124
rect -1964 8090 -1930 8124
rect -1896 8090 -1862 8124
rect -1828 8090 -1794 8124
rect -1760 8090 -1726 8124
rect -1692 8090 -1658 8124
rect -1624 8090 -1590 8124
rect -1556 8090 -1522 8124
rect -1488 8090 -1454 8124
rect -1420 8090 -1386 8124
rect -1352 8090 -1318 8124
rect -1284 8090 -1250 8124
rect -1216 8090 -1182 8124
rect -1148 8090 -1114 8124
rect -1080 8090 -1046 8124
rect -1012 8090 -978 8124
rect -944 8090 -910 8124
rect -876 8090 -842 8124
rect -808 8090 -774 8124
rect -740 8090 -706 8124
rect -672 8090 -638 8124
rect -604 8090 -570 8124
rect -536 8090 -502 8124
rect -468 8090 -434 8124
rect -400 8090 -366 8124
rect -332 8090 -298 8124
rect -264 8090 -230 8124
rect -196 8090 -162 8124
rect -128 8090 -94 8124
rect -60 8090 -26 8124
rect 8 8090 42 8124
rect 76 8090 110 8124
rect 144 8090 178 8124
rect 212 8090 246 8124
rect 280 8090 314 8124
rect 348 8090 382 8124
rect 416 8090 450 8124
rect 484 8090 518 8124
rect 552 8090 586 8124
rect 620 8090 654 8124
rect 688 8090 722 8124
rect 756 8090 790 8124
rect 824 8090 858 8124
rect 892 8090 926 8124
rect 960 8090 994 8124
rect 1028 8090 1062 8124
rect 1096 8090 1142 8124
rect 1176 8090 1210 8124
rect 1244 8090 1278 8124
rect 1312 8090 1346 8124
rect 1380 8090 1414 8124
rect 1448 8090 1552 8124
rect -2322 8002 -2288 8090
rect -2322 7934 -2288 7968
rect 1518 8002 1552 8090
rect -2322 7866 -2288 7900
rect -2322 7798 -2288 7832
rect -2322 7730 -2288 7764
rect 1518 7934 1552 7968
rect 1518 7866 1552 7900
rect 1518 7798 1552 7832
rect -2322 7662 -2288 7696
rect 1518 7730 1552 7764
rect 1518 7662 1552 7696
rect -2322 7594 -2288 7628
rect -2322 7526 -2288 7560
rect 1518 7594 1552 7628
rect -2322 7458 -2288 7492
rect -2322 7390 -2288 7424
rect -2322 7322 -2288 7356
rect 1518 7526 1552 7560
rect 1518 7458 1552 7492
rect 9741 7603 10350 7761
rect 9741 7501 9914 7603
rect 10288 7501 10350 7603
rect 1518 7390 1552 7424
rect -2322 7254 -2288 7288
rect 1518 7322 1552 7356
rect 1518 7254 1552 7288
rect -2322 7186 -2288 7220
rect -2322 7118 -2288 7152
rect 1518 7186 1552 7220
rect 1518 7118 1552 7152
rect -2322 7050 -2288 7084
rect -2322 6982 -2288 7016
rect -2322 6914 -2288 6948
rect 1518 7050 1552 7084
rect 1518 6982 1552 7016
rect 1518 6914 1552 6948
rect -2322 6846 -2288 6880
rect 1518 6846 1552 6880
rect -2322 6778 -2288 6812
rect -2322 6710 -2288 6744
rect 1518 6778 1552 6812
rect 1518 6710 1552 6744
rect -2322 6642 -2288 6676
rect -2322 6574 -2288 6608
rect -2322 6506 -2288 6540
rect 1518 6642 1552 6676
rect 1518 6574 1552 6608
rect 1518 6506 1552 6540
rect -2322 6438 -2288 6472
rect 1518 6438 1552 6472
rect -2322 6370 -2288 6404
rect 1518 6370 1552 6404
rect -2322 6302 -2288 6336
rect 1518 6302 1552 6336
rect -2322 6234 -2288 6268
rect -2322 6166 -2288 6200
rect -2322 6098 -2288 6132
rect 1518 6234 1552 6268
rect 1518 6166 1552 6200
rect 1518 6098 1552 6132
rect -2322 6030 -2288 6064
rect -2322 5962 -2288 5996
rect 1518 6030 1552 6064
rect 1518 5962 1552 5996
rect -2322 5894 -2288 5928
rect 1518 5894 1552 5928
rect -2322 5826 -2288 5860
rect -2322 5758 -2288 5792
rect -2322 5690 -2288 5724
rect 1518 5826 1552 5860
rect 1518 5758 1552 5792
rect 1518 5690 1552 5724
rect -2322 5622 -2288 5656
rect -2322 5554 -2288 5588
rect 1518 5622 1552 5656
rect 1518 5554 1552 5588
rect -2322 5486 -2288 5520
rect -2322 5418 -2288 5452
rect 1518 5486 1552 5520
rect -2322 5350 -2288 5384
rect -2322 5282 -2288 5316
rect -2322 5214 -2288 5248
rect 1518 5418 1552 5452
rect 1518 5350 1552 5384
rect 1518 5282 1552 5316
rect -2322 5146 -2288 5180
rect 1518 5214 1552 5248
rect 1518 5146 1552 5180
rect -2322 5078 -2288 5112
rect -2322 5010 -2288 5044
rect 1518 5078 1552 5112
rect -2322 4942 -2288 4976
rect -2322 4874 -2288 4908
rect -2322 4806 -2288 4840
rect 1518 5010 1552 5044
rect 1518 4942 1552 4976
rect 1518 4874 1552 4908
rect -2322 4738 -2288 4772
rect 1518 4806 1552 4840
rect 1518 4738 1552 4772
rect -2322 4670 -2288 4704
rect -2322 4602 -2288 4636
rect 1518 4670 1552 4704
rect -2322 4534 -2288 4568
rect -2322 4466 -2288 4500
rect -2322 4398 -2288 4432
rect 1518 4602 1552 4636
rect 1518 4534 1552 4568
rect 1518 4466 1552 4500
rect -2322 4330 -2288 4364
rect 1518 4398 1552 4432
rect 1518 4330 1552 4364
rect -2322 4262 -2288 4296
rect -2322 4194 -2288 4228
rect 1518 4262 1552 4296
rect 1518 4194 1552 4228
rect -2322 4126 -2288 4160
rect -2322 4058 -2288 4092
rect -2322 3990 -2288 4024
rect 1518 4126 1552 4160
rect 1518 4058 1552 4092
rect 1518 3990 1552 4024
rect 3508 7451 3628 7485
rect 3662 7451 3696 7485
rect 3730 7451 3764 7485
rect 3798 7451 3832 7485
rect 3866 7451 3900 7485
rect 3934 7451 3968 7485
rect 4002 7451 4036 7485
rect 4070 7451 4104 7485
rect 4138 7451 4172 7485
rect 4206 7451 4240 7485
rect 4274 7451 4308 7485
rect 4342 7451 4376 7485
rect 4410 7451 4444 7485
rect 4478 7451 4512 7485
rect 4546 7451 4580 7485
rect 4614 7451 4648 7485
rect 4682 7451 4716 7485
rect 4750 7451 4784 7485
rect 4818 7451 4852 7485
rect 4886 7451 4920 7485
rect 4954 7451 4988 7485
rect 5022 7451 5056 7485
rect 5090 7451 5124 7485
rect 5158 7451 5192 7485
rect 5226 7451 5260 7485
rect 5294 7451 5328 7485
rect 5362 7451 5396 7485
rect 5430 7451 5464 7485
rect 5498 7451 5532 7485
rect 5566 7451 5600 7485
rect 5634 7451 5668 7485
rect 5702 7451 5736 7485
rect 5770 7451 5804 7485
rect 5838 7451 5872 7485
rect 5906 7451 5940 7485
rect 5974 7451 6008 7485
rect 6042 7451 6076 7485
rect 6110 7451 6144 7485
rect 6178 7451 6212 7485
rect 6246 7451 6350 7485
rect 3508 7363 3542 7451
rect 3508 7295 3542 7329
rect 6316 7363 6350 7451
rect 9741 7364 10350 7501
rect 3508 7227 3542 7261
rect 3508 7159 3542 7193
rect 3508 7091 3542 7125
rect 6316 7295 6350 7329
rect 6316 7227 6350 7261
rect 6316 7159 6350 7193
rect 3508 7023 3542 7057
rect 6316 7091 6350 7125
rect 6316 7023 6350 7057
rect 3508 6955 3542 6989
rect 3508 6887 3542 6921
rect 6316 6955 6350 6989
rect 3508 6819 3542 6853
rect 3508 6751 3542 6785
rect 3508 6683 3542 6717
rect 6316 6887 6350 6921
rect 6316 6819 6350 6853
rect 6316 6751 6350 6785
rect 3508 6615 3542 6649
rect 6316 6683 6350 6717
rect 6316 6615 6350 6649
rect 3508 6547 3542 6581
rect 3508 6479 3542 6513
rect 6316 6479 6350 6581
rect 3508 6411 3542 6445
rect 3508 6343 3542 6377
rect 3508 6275 3542 6309
rect 6316 6411 6350 6445
rect 6316 6343 6350 6377
rect 6316 6275 6350 6309
rect 3508 6207 3542 6241
rect 6316 6207 6350 6241
rect 3508 6139 3542 6173
rect 3508 6071 3542 6105
rect 6316 6139 6350 6173
rect 6316 6071 6350 6105
rect 3508 6003 3542 6037
rect 3508 5935 3542 5969
rect 3508 5867 3542 5901
rect 6316 6003 6350 6037
rect 6316 5935 6350 5969
rect 6316 5867 6350 5901
rect 3508 5799 3542 5833
rect 6316 5799 6350 5833
rect 3508 5731 3542 5765
rect 6316 5731 6350 5765
rect 3508 5663 3542 5697
rect 6316 5663 6350 5697
rect 3508 5595 3542 5629
rect 3508 5527 3542 5561
rect 3508 5459 3542 5493
rect 6316 5595 6350 5629
rect 6316 5527 6350 5561
rect 6316 5459 6350 5493
rect 3508 5391 3542 5425
rect 3508 5323 3542 5357
rect 6316 5391 6350 5425
rect 6316 5323 6350 5357
rect 3508 5255 3542 5289
rect 6316 5255 6350 5289
rect 3508 5187 3542 5221
rect 3508 5119 3542 5153
rect 3508 5051 3542 5085
rect 6316 5187 6350 5221
rect 6316 5119 6350 5153
rect 6316 5051 6350 5085
rect 3508 4983 3542 5017
rect 3508 4915 3542 4949
rect 6316 4915 6350 5017
rect 3508 4847 3542 4881
rect 3508 4779 3542 4813
rect 6316 4847 6350 4881
rect 3508 4711 3542 4745
rect 3508 4643 3542 4677
rect 3508 4575 3542 4609
rect 6316 4779 6350 4813
rect 6316 4711 6350 4745
rect 6316 4643 6350 4677
rect 3508 4507 3542 4541
rect 6316 4575 6350 4609
rect 6316 4507 6350 4541
rect 3508 4439 3542 4473
rect 3508 4371 3542 4405
rect 6316 4439 6350 4473
rect 3508 4303 3542 4337
rect 3508 4235 3542 4269
rect 3508 4167 3542 4201
rect 6316 4371 6350 4405
rect 6316 4303 6350 4337
rect 6316 4235 6350 4269
rect 3508 4045 3542 4133
rect 6316 4167 6350 4201
rect 6316 4045 6350 4133
rect 3508 4011 3628 4045
rect 3662 4011 3696 4045
rect 3730 4011 3764 4045
rect 3798 4011 3832 4045
rect 3866 4011 3900 4045
rect 3934 4011 3968 4045
rect 4002 4011 4036 4045
rect 4070 4011 4104 4045
rect 4138 4011 4172 4045
rect 4206 4011 4240 4045
rect 4274 4011 4308 4045
rect 4342 4011 4376 4045
rect 4410 4011 4444 4045
rect 4478 4011 4512 4045
rect 4546 4011 4580 4045
rect 4614 4011 4648 4045
rect 4682 4011 4716 4045
rect 4750 4011 4784 4045
rect 4818 4011 4852 4045
rect 4886 4011 4920 4045
rect 4954 4011 4988 4045
rect 5022 4011 5056 4045
rect 5090 4011 5124 4045
rect 5158 4011 5192 4045
rect 5226 4011 5260 4045
rect 5294 4011 5328 4045
rect 5362 4011 5396 4045
rect 5430 4011 5464 4045
rect 5498 4011 5532 4045
rect 5566 4011 5600 4045
rect 5634 4011 5668 4045
rect 5702 4011 5736 4045
rect 5770 4011 5804 4045
rect 5838 4011 5872 4045
rect 5906 4011 5940 4045
rect 5974 4011 6008 4045
rect 6042 4011 6076 4045
rect 6110 4011 6144 4045
rect 6178 4011 6212 4045
rect 6246 4011 6350 4045
rect 8244 7040 8364 7074
rect 8398 7040 8432 7074
rect 8466 7040 8500 7074
rect 8534 7040 8568 7074
rect 8602 7040 8636 7074
rect 8670 7040 8704 7074
rect 8738 7040 8772 7074
rect 8806 7040 8840 7074
rect 8874 7040 8908 7074
rect 8942 7040 8976 7074
rect 9010 7040 9044 7074
rect 9078 7040 9112 7074
rect 9146 7040 9180 7074
rect 9214 7040 9248 7074
rect 9282 7040 9316 7074
rect 9350 7040 9384 7074
rect 9418 7040 9452 7074
rect 9486 7040 9520 7074
rect 9554 7040 9588 7074
rect 9622 7040 9656 7074
rect 9690 7040 9724 7074
rect 9758 7040 9792 7074
rect 9826 7040 9860 7074
rect 9894 7040 9928 7074
rect 9962 7040 10054 7074
rect 8244 6952 8278 7040
rect 8244 6884 8278 6918
rect 10020 6952 10054 7040
rect 8244 6816 8278 6850
rect 8244 6748 8278 6782
rect 8244 6680 8278 6714
rect 10020 6884 10054 6918
rect 10020 6816 10054 6850
rect 10020 6748 10054 6782
rect 8244 6612 8278 6646
rect 10020 6680 10054 6714
rect 10020 6612 10054 6646
rect 8244 6544 8278 6578
rect 8244 6476 8278 6510
rect 10020 6544 10054 6578
rect 8244 6408 8278 6442
rect 8244 6340 8278 6374
rect 8244 6272 8278 6306
rect 10020 6476 10054 6510
rect 10020 6408 10054 6442
rect 10020 6340 10054 6374
rect 8244 6204 8278 6238
rect 10020 6272 10054 6306
rect 10020 6204 10054 6238
rect 8244 6136 8278 6170
rect 8244 6068 8278 6102
rect 10020 6068 10054 6170
rect 8244 6000 8278 6034
rect 8244 5932 8278 5966
rect 8244 5864 8278 5898
rect 10020 6000 10054 6034
rect 10020 5932 10054 5966
rect 10020 5864 10054 5898
rect 8244 5796 8278 5830
rect 10020 5796 10054 5830
rect 8244 5728 8278 5762
rect 8244 5660 8278 5694
rect 10020 5728 10054 5762
rect 10020 5660 10054 5694
rect 8244 5592 8278 5626
rect 8244 5524 8278 5558
rect 8244 5456 8278 5490
rect 10020 5592 10054 5626
rect 10020 5524 10054 5558
rect 10020 5456 10054 5490
rect 8244 5388 8278 5422
rect 10020 5388 10054 5422
rect 8244 5320 8278 5354
rect 10020 5320 10054 5354
rect 8244 5252 8278 5286
rect 10020 5252 10054 5286
rect 8244 5184 8278 5218
rect 8244 5116 8278 5150
rect 8244 5048 8278 5082
rect 10020 5184 10054 5218
rect 10020 5116 10054 5150
rect 10020 5048 10054 5082
rect 8244 4980 8278 5014
rect 8244 4912 8278 4946
rect 10020 4980 10054 5014
rect 10020 4912 10054 4946
rect 8244 4844 8278 4878
rect 10020 4844 10054 4878
rect 8244 4776 8278 4810
rect 8244 4708 8278 4742
rect 8244 4640 8278 4674
rect 10020 4776 10054 4810
rect 10020 4708 10054 4742
rect 10020 4640 10054 4674
rect 8244 4572 8278 4606
rect 8244 4504 8278 4538
rect 10020 4504 10054 4606
rect 8244 4436 8278 4470
rect 8244 4368 8278 4402
rect 10020 4436 10054 4470
rect 8244 4300 8278 4334
rect 8244 4232 8278 4266
rect 8244 4164 8278 4198
rect 10020 4368 10054 4402
rect 10020 4300 10054 4334
rect 10020 4232 10054 4266
rect 8244 4052 8278 4130
rect 10020 4164 10054 4198
rect 10020 4052 10054 4130
rect 8244 4018 8364 4052
rect 8398 4018 8432 4052
rect 8466 4018 8500 4052
rect 8534 4018 8568 4052
rect 8602 4018 8636 4052
rect 8670 4018 8704 4052
rect 8738 4018 8772 4052
rect 8806 4018 8840 4052
rect 8874 4018 8908 4052
rect 8942 4018 8976 4052
rect 9010 4018 9044 4052
rect 9078 4018 9112 4052
rect 9146 4018 9180 4052
rect 9214 4018 9248 4052
rect 9282 4018 9316 4052
rect 9350 4018 9384 4052
rect 9418 4018 9452 4052
rect 9486 4018 9520 4052
rect 9554 4018 9588 4052
rect 9622 4018 9656 4052
rect 9690 4018 9724 4052
rect 9758 4018 9792 4052
rect 9826 4018 9860 4052
rect 9894 4018 10054 4052
rect -2322 3848 -2288 3956
rect 1518 3848 1552 3956
rect -2322 3814 -2202 3848
rect -2168 3814 -2134 3848
rect -2100 3814 -2066 3848
rect -2032 3814 -1998 3848
rect -1964 3814 -1930 3848
rect -1896 3814 -1862 3848
rect -1828 3814 -1794 3848
rect -1760 3814 -1726 3848
rect -1692 3814 -1658 3848
rect -1624 3814 -1590 3848
rect -1556 3814 -1522 3848
rect -1488 3814 -1454 3848
rect -1420 3814 -1386 3848
rect -1352 3814 -1318 3848
rect -1284 3814 -1250 3848
rect -1216 3814 -1182 3848
rect -1148 3814 -1114 3848
rect -1080 3814 -1046 3848
rect -1012 3814 -978 3848
rect -944 3814 -910 3848
rect -876 3814 -842 3848
rect -808 3814 -774 3848
rect -740 3814 -706 3848
rect -672 3814 -638 3848
rect -604 3814 -570 3848
rect -536 3814 -502 3848
rect -468 3814 -434 3848
rect -400 3814 -366 3848
rect -332 3814 -298 3848
rect -264 3814 -230 3848
rect -196 3814 -162 3848
rect -128 3814 -94 3848
rect -60 3814 -26 3848
rect 8 3814 42 3848
rect 76 3814 110 3848
rect 144 3814 178 3848
rect 212 3814 246 3848
rect 280 3814 314 3848
rect 348 3814 382 3848
rect 416 3814 450 3848
rect 484 3814 518 3848
rect 552 3814 586 3848
rect 620 3814 654 3848
rect 688 3814 722 3848
rect 756 3814 790 3848
rect 824 3814 858 3848
rect 892 3814 926 3848
rect 960 3814 994 3848
rect 1028 3814 1062 3848
rect 1096 3814 1130 3848
rect 1164 3814 1198 3848
rect 1232 3814 1266 3848
rect 1300 3814 1334 3848
rect 1368 3814 1402 3848
rect 1436 3814 1552 3848
<< nsubdiff >>
rect 6895 10947 7015 10981
rect 7049 10947 7083 10981
rect 7117 10947 7151 10981
rect 7185 10947 7219 10981
rect 7253 10947 7287 10981
rect 7321 10947 7355 10981
rect 7389 10947 7423 10981
rect 7457 10947 7491 10981
rect 7525 10947 7559 10981
rect 7593 10947 7627 10981
rect 7661 10947 7695 10981
rect 7729 10947 7763 10981
rect 7797 10947 7831 10981
rect 7865 10947 7899 10981
rect 7933 10947 7967 10981
rect 8001 10947 8035 10981
rect 8069 10947 8103 10981
rect 8137 10947 8171 10981
rect 8205 10947 8239 10981
rect 8273 10947 8307 10981
rect 8341 10947 8375 10981
rect 8409 10947 8443 10981
rect 8477 10947 8511 10981
rect 8545 10947 8579 10981
rect 8613 10947 8705 10981
rect -1353 10629 -1233 10663
rect -1199 10629 -1165 10663
rect -1131 10629 -1097 10663
rect -1063 10629 -1029 10663
rect -995 10629 -961 10663
rect -927 10629 -893 10663
rect -859 10629 -825 10663
rect -791 10629 -757 10663
rect -723 10629 -689 10663
rect -655 10629 -621 10663
rect -587 10629 -553 10663
rect -519 10629 -485 10663
rect -451 10629 -417 10663
rect -383 10629 -349 10663
rect -315 10629 -281 10663
rect -247 10629 -213 10663
rect -179 10629 -145 10663
rect -111 10629 -77 10663
rect -43 10629 -9 10663
rect 25 10629 59 10663
rect 93 10629 127 10663
rect 161 10629 195 10663
rect 229 10629 263 10663
rect 297 10629 331 10663
rect 365 10629 457 10663
rect -1353 10551 -1319 10629
rect -1353 10483 -1319 10517
rect 423 10551 457 10629
rect 423 10483 457 10517
rect -1353 10415 -1319 10449
rect -1353 10347 -1319 10381
rect -1353 10279 -1319 10313
rect 423 10415 457 10449
rect 423 10347 457 10381
rect -1353 10211 -1319 10245
rect 423 10279 457 10313
rect 423 10211 457 10245
rect -1353 10143 -1319 10177
rect 423 10143 457 10177
rect -1353 10075 -1319 10109
rect 423 10075 457 10109
rect -1353 10007 -1319 10041
rect -1353 9939 -1319 9973
rect -1353 9871 -1319 9905
rect 423 10007 457 10041
rect 423 9939 457 9973
rect 423 9871 457 9905
rect -1353 9803 -1319 9837
rect -1353 9735 -1319 9769
rect 423 9803 457 9837
rect 423 9735 457 9769
rect -1353 9667 -1319 9701
rect -1353 9599 -1319 9633
rect 423 9667 457 9701
rect -1353 9531 -1319 9565
rect -1353 9463 -1319 9497
rect -1353 9395 -1319 9429
rect 423 9599 457 9633
rect 423 9531 457 9565
rect 423 9463 457 9497
rect -1353 9327 -1319 9361
rect 423 9395 457 9429
rect 423 9327 457 9361
rect -1353 9259 -1319 9293
rect -1353 9191 -1319 9225
rect 423 9259 457 9293
rect 423 9191 457 9225
rect -1353 9123 -1319 9157
rect -1353 9055 -1319 9089
rect -1353 8987 -1319 9021
rect 423 9123 457 9157
rect 423 9055 457 9089
rect 423 8987 457 9021
rect -1353 8919 -1319 8953
rect -1353 8823 -1319 8885
rect 423 8919 457 8953
rect 423 8823 457 8885
rect -1353 8789 -1233 8823
rect -1199 8789 -1165 8823
rect -1131 8789 -1097 8823
rect -1063 8789 -1029 8823
rect -995 8789 -961 8823
rect -927 8789 -893 8823
rect -859 8789 -825 8823
rect -791 8789 -757 8823
rect -723 8789 -689 8823
rect -655 8789 -621 8823
rect -587 8789 -553 8823
rect -519 8789 -485 8823
rect -451 8789 -417 8823
rect -383 8789 -349 8823
rect -315 8789 -281 8823
rect -247 8789 -213 8823
rect -179 8789 -145 8823
rect -111 8789 -77 8823
rect -43 8789 -9 8823
rect 25 8789 59 8823
rect 93 8789 127 8823
rect 161 8789 195 8823
rect 229 8789 263 8823
rect 297 8789 331 8823
rect 365 8789 457 8823
rect 6895 10869 6929 10947
rect 6895 10801 6929 10835
rect 8671 10869 8705 10947
rect 8671 10801 8705 10835
rect 6895 10733 6929 10767
rect 6895 10665 6929 10699
rect 6895 10597 6929 10631
rect 8671 10733 8705 10767
rect 8671 10665 8705 10699
rect 6895 10529 6929 10563
rect 8671 10597 8705 10631
rect 8671 10529 8705 10563
rect 6895 10461 6929 10495
rect 8671 10461 8705 10495
rect 6895 10393 6929 10427
rect 8671 10393 8705 10427
rect 6895 10325 6929 10359
rect 6895 10257 6929 10291
rect 6895 10189 6929 10223
rect 8671 10325 8705 10359
rect 8671 10257 8705 10291
rect 8671 10189 8705 10223
rect 6895 10121 6929 10155
rect 6895 10053 6929 10087
rect 8671 10121 8705 10155
rect 8671 10053 8705 10087
rect 6895 9985 6929 10019
rect 6895 9917 6929 9951
rect 8671 9985 8705 10019
rect 6895 9849 6929 9883
rect 6895 9781 6929 9815
rect 6895 9713 6929 9747
rect 8671 9917 8705 9951
rect 8671 9849 8705 9883
rect 8671 9781 8705 9815
rect 6895 9645 6929 9679
rect 8671 9713 8705 9747
rect 8671 9645 8705 9679
rect 6895 9577 6929 9611
rect 6895 9509 6929 9543
rect 8671 9577 8705 9611
rect 8671 9509 8705 9543
rect 6895 9441 6929 9475
rect 6895 9373 6929 9407
rect 6895 9305 6929 9339
rect 8671 9441 8705 9475
rect 8671 9373 8705 9407
rect 8671 9305 8705 9339
rect 6895 9237 6929 9271
rect 6895 9169 6929 9203
rect 8671 9237 8705 9271
rect 8671 9169 8705 9203
rect 6895 9101 6929 9135
rect 6895 9033 6929 9067
rect 8671 9101 8705 9135
rect 6895 8965 6929 8999
rect 6895 8897 6929 8931
rect 6895 8829 6929 8863
rect 8671 9033 8705 9067
rect 8671 8965 8705 8999
rect 8671 8897 8705 8931
rect 6895 8761 6929 8795
rect 8671 8829 8705 8863
rect 8671 8761 8705 8795
rect 6895 8693 6929 8727
rect 6895 8625 6929 8659
rect 8671 8693 8705 8727
rect 8671 8625 8705 8659
rect 6895 8557 6929 8591
rect 6895 8489 6929 8523
rect 6895 8421 6929 8455
rect 8671 8557 8705 8591
rect 8671 8489 8705 8523
rect 8671 8421 8705 8455
rect 6895 8353 6929 8387
rect 8671 8353 8705 8387
rect 6895 8285 6929 8319
rect 8671 8285 8705 8319
rect 6895 8217 6929 8251
rect 6895 8149 6929 8183
rect 8671 8217 8705 8251
rect 6895 8081 6929 8115
rect 6895 8013 6929 8047
rect 8671 8149 8705 8183
rect 8671 8081 8705 8115
rect 8671 8013 8705 8047
rect 6895 7945 6929 7979
rect 6895 7833 6929 7911
rect 8671 7945 8705 7979
rect 8671 7833 8705 7911
rect 6895 7799 7015 7833
rect 7049 7799 7083 7833
rect 7117 7799 7151 7833
rect 7185 7799 7219 7833
rect 7253 7799 7287 7833
rect 7321 7799 7355 7833
rect 7389 7799 7423 7833
rect 7457 7799 7491 7833
rect 7525 7799 7559 7833
rect 7593 7799 7627 7833
rect 7661 7799 7695 7833
rect 7729 7799 7763 7833
rect 7797 7799 7831 7833
rect 7865 7799 7899 7833
rect 7933 7799 7967 7833
rect 8001 7799 8035 7833
rect 8069 7799 8103 7833
rect 8137 7799 8171 7833
rect 8205 7799 8239 7833
rect 8273 7799 8307 7833
rect 8341 7799 8375 7833
rect 8409 7799 8443 7833
rect 8477 7799 8511 7833
rect 8545 7799 8579 7833
rect 8613 7799 8705 7833
<< psubdiffcont >>
rect 3089 10839 3123 10873
rect 3157 10839 3191 10873
rect 3225 10839 3259 10873
rect 3293 10839 3327 10873
rect 3361 10839 3395 10873
rect 3429 10839 3463 10873
rect 3497 10839 3531 10873
rect 3565 10839 3599 10873
rect 3633 10839 3667 10873
rect 3701 10839 3735 10873
rect 3769 10839 3803 10873
rect 3837 10839 3871 10873
rect 3905 10839 3939 10873
rect 3973 10839 4007 10873
rect 4041 10839 4075 10873
rect 4109 10839 4143 10873
rect 4177 10839 4211 10873
rect 4245 10839 4279 10873
rect 4313 10839 4347 10873
rect 4381 10839 4415 10873
rect 4449 10839 4483 10873
rect 4517 10839 4551 10873
rect 4585 10839 4619 10873
rect 4653 10839 4687 10873
rect 4721 10839 4755 10873
rect 4789 10839 4823 10873
rect 4857 10839 4891 10873
rect 4925 10839 4959 10873
rect 4993 10839 5027 10873
rect 5061 10839 5095 10873
rect 5129 10839 5163 10873
rect 2969 10737 3003 10771
rect 2969 10669 3003 10703
rect 5262 10737 5296 10771
rect 2969 10601 3003 10635
rect 2969 10533 3003 10567
rect 5262 10669 5296 10703
rect 5262 10601 5296 10635
rect 5262 10533 5296 10567
rect 2969 10465 3003 10499
rect 2969 10397 3003 10431
rect 5262 10465 5296 10499
rect 5262 10397 5296 10431
rect 2969 10329 3003 10363
rect 2969 10261 3003 10295
rect 5262 10329 5296 10363
rect 2969 10193 3003 10227
rect 2969 10125 3003 10159
rect 2969 10057 3003 10091
rect 5262 10261 5296 10295
rect 5262 10193 5296 10227
rect 5262 10125 5296 10159
rect 2969 9989 3003 10023
rect 5262 10057 5296 10091
rect 2969 9921 3003 9955
rect 5262 9989 5296 10023
rect 2969 9853 3003 9887
rect 5262 9921 5296 9955
rect 2969 9785 3003 9819
rect 2969 9717 3003 9751
rect 2969 9649 3003 9683
rect 5262 9853 5296 9887
rect 5262 9785 5296 9819
rect 5262 9717 5296 9751
rect 2969 9581 3003 9615
rect 5262 9649 5296 9683
rect 5262 9581 5296 9615
rect 2969 9513 3003 9547
rect 2969 9445 3003 9479
rect 5262 9513 5296 9547
rect 5262 9445 5296 9479
rect 2969 9377 3003 9411
rect 2969 9309 3003 9343
rect 2969 9241 3003 9275
rect 5262 9377 5296 9411
rect 5262 9309 5296 9343
rect 2969 9173 3003 9207
rect 5262 9241 5296 9275
rect 5262 9173 5296 9207
rect 2969 9105 3003 9139
rect 2969 9037 3003 9071
rect 5262 9105 5296 9139
rect 5262 9037 5296 9071
rect 2969 8969 3003 9003
rect 2969 8901 3003 8935
rect 2969 8833 3003 8867
rect 5262 8969 5296 9003
rect 5262 8901 5296 8935
rect 5262 8833 5296 8867
rect 2969 8765 3003 8799
rect 5262 8765 5296 8799
rect 2969 8697 3003 8731
rect 5262 8697 5296 8731
rect 2969 8629 3003 8663
rect 5262 8629 5296 8663
rect 2969 8561 3003 8595
rect 2969 8493 3003 8527
rect 2969 8425 3003 8459
rect 5262 8561 5296 8595
rect 5262 8493 5296 8527
rect 5262 8425 5296 8459
rect 2969 8357 3003 8391
rect 5262 8357 5296 8391
rect 3089 8234 3123 8268
rect 3157 8234 3191 8268
rect 3225 8234 3259 8268
rect 3293 8234 3327 8268
rect 3361 8234 3395 8268
rect 3429 8234 3463 8268
rect 3497 8234 3531 8268
rect 3565 8234 3599 8268
rect 3633 8234 3667 8268
rect 3701 8234 3735 8268
rect 3769 8234 3803 8268
rect 3837 8234 3871 8268
rect 3905 8234 3939 8268
rect 3973 8234 4007 8268
rect 4041 8234 4075 8268
rect 4109 8234 4143 8268
rect 4177 8234 4211 8268
rect 4245 8234 4279 8268
rect 4313 8234 4347 8268
rect 4381 8234 4415 8268
rect 4449 8234 4483 8268
rect 4517 8234 4551 8268
rect 4585 8234 4619 8268
rect 4653 8234 4687 8268
rect 4721 8234 4755 8268
rect 4789 8234 4823 8268
rect 4857 8234 4891 8268
rect 4925 8234 4959 8268
rect 4993 8234 5027 8268
rect 5061 8234 5095 8268
rect 5129 8234 5163 8268
rect -2202 8090 -2168 8124
rect -2134 8090 -2100 8124
rect -2066 8090 -2032 8124
rect -1998 8090 -1964 8124
rect -1930 8090 -1896 8124
rect -1862 8090 -1828 8124
rect -1794 8090 -1760 8124
rect -1726 8090 -1692 8124
rect -1658 8090 -1624 8124
rect -1590 8090 -1556 8124
rect -1522 8090 -1488 8124
rect -1454 8090 -1420 8124
rect -1386 8090 -1352 8124
rect -1318 8090 -1284 8124
rect -1250 8090 -1216 8124
rect -1182 8090 -1148 8124
rect -1114 8090 -1080 8124
rect -1046 8090 -1012 8124
rect -978 8090 -944 8124
rect -910 8090 -876 8124
rect -842 8090 -808 8124
rect -774 8090 -740 8124
rect -706 8090 -672 8124
rect -638 8090 -604 8124
rect -570 8090 -536 8124
rect -502 8090 -468 8124
rect -434 8090 -400 8124
rect -366 8090 -332 8124
rect -298 8090 -264 8124
rect -230 8090 -196 8124
rect -162 8090 -128 8124
rect -94 8090 -60 8124
rect -26 8090 8 8124
rect 42 8090 76 8124
rect 110 8090 144 8124
rect 178 8090 212 8124
rect 246 8090 280 8124
rect 314 8090 348 8124
rect 382 8090 416 8124
rect 450 8090 484 8124
rect 518 8090 552 8124
rect 586 8090 620 8124
rect 654 8090 688 8124
rect 722 8090 756 8124
rect 790 8090 824 8124
rect 858 8090 892 8124
rect 926 8090 960 8124
rect 994 8090 1028 8124
rect 1062 8090 1096 8124
rect 1142 8090 1176 8124
rect 1210 8090 1244 8124
rect 1278 8090 1312 8124
rect 1346 8090 1380 8124
rect 1414 8090 1448 8124
rect -2322 7968 -2288 8002
rect 1518 7968 1552 8002
rect -2322 7900 -2288 7934
rect -2322 7832 -2288 7866
rect -2322 7764 -2288 7798
rect 1518 7900 1552 7934
rect 1518 7832 1552 7866
rect 1518 7764 1552 7798
rect -2322 7696 -2288 7730
rect 1518 7696 1552 7730
rect -2322 7628 -2288 7662
rect 1518 7628 1552 7662
rect -2322 7560 -2288 7594
rect 1518 7560 1552 7594
rect -2322 7492 -2288 7526
rect -2322 7424 -2288 7458
rect -2322 7356 -2288 7390
rect 1518 7492 1552 7526
rect 9914 7501 10288 7603
rect 1518 7424 1552 7458
rect 1518 7356 1552 7390
rect -2322 7288 -2288 7322
rect -2322 7220 -2288 7254
rect 1518 7288 1552 7322
rect 1518 7220 1552 7254
rect -2322 7152 -2288 7186
rect -2322 7084 -2288 7118
rect 1518 7152 1552 7186
rect -2322 7016 -2288 7050
rect -2322 6948 -2288 6982
rect 1518 7084 1552 7118
rect 1518 7016 1552 7050
rect 1518 6948 1552 6982
rect -2322 6880 -2288 6914
rect -2322 6812 -2288 6846
rect 1518 6880 1552 6914
rect 1518 6812 1552 6846
rect -2322 6744 -2288 6778
rect -2322 6676 -2288 6710
rect 1518 6744 1552 6778
rect -2322 6608 -2288 6642
rect -2322 6540 -2288 6574
rect -2322 6472 -2288 6506
rect 1518 6676 1552 6710
rect 1518 6608 1552 6642
rect 1518 6540 1552 6574
rect -2322 6404 -2288 6438
rect 1518 6472 1552 6506
rect -2322 6336 -2288 6370
rect 1518 6404 1552 6438
rect -2322 6268 -2288 6302
rect 1518 6336 1552 6370
rect -2322 6200 -2288 6234
rect -2322 6132 -2288 6166
rect -2322 6064 -2288 6098
rect 1518 6268 1552 6302
rect 1518 6200 1552 6234
rect 1518 6132 1552 6166
rect -2322 5996 -2288 6030
rect 1518 6064 1552 6098
rect 1518 5996 1552 6030
rect -2322 5928 -2288 5962
rect -2322 5860 -2288 5894
rect 1518 5928 1552 5962
rect 1518 5860 1552 5894
rect -2322 5792 -2288 5826
rect -2322 5724 -2288 5758
rect -2322 5656 -2288 5690
rect 1518 5792 1552 5826
rect 1518 5724 1552 5758
rect -2322 5588 -2288 5622
rect 1518 5656 1552 5690
rect 1518 5588 1552 5622
rect -2322 5520 -2288 5554
rect -2322 5452 -2288 5486
rect 1518 5520 1552 5554
rect 1518 5452 1552 5486
rect -2322 5384 -2288 5418
rect -2322 5316 -2288 5350
rect -2322 5248 -2288 5282
rect 1518 5384 1552 5418
rect 1518 5316 1552 5350
rect 1518 5248 1552 5282
rect -2322 5180 -2288 5214
rect 1518 5180 1552 5214
rect -2322 5112 -2288 5146
rect 1518 5112 1552 5146
rect -2322 5044 -2288 5078
rect 1518 5044 1552 5078
rect -2322 4976 -2288 5010
rect -2322 4908 -2288 4942
rect -2322 4840 -2288 4874
rect 1518 4976 1552 5010
rect 1518 4908 1552 4942
rect 1518 4840 1552 4874
rect -2322 4772 -2288 4806
rect -2322 4704 -2288 4738
rect 1518 4772 1552 4806
rect 1518 4704 1552 4738
rect -2322 4636 -2288 4670
rect 1518 4636 1552 4670
rect -2322 4568 -2288 4602
rect -2322 4500 -2288 4534
rect -2322 4432 -2288 4466
rect 1518 4568 1552 4602
rect 1518 4500 1552 4534
rect 1518 4432 1552 4466
rect -2322 4364 -2288 4398
rect -2322 4296 -2288 4330
rect 1518 4364 1552 4398
rect 1518 4296 1552 4330
rect -2322 4228 -2288 4262
rect -2322 4160 -2288 4194
rect 1518 4228 1552 4262
rect -2322 4092 -2288 4126
rect -2322 4024 -2288 4058
rect -2322 3956 -2288 3990
rect 1518 4160 1552 4194
rect 1518 4092 1552 4126
rect 1518 4024 1552 4058
rect 3628 7451 3662 7485
rect 3696 7451 3730 7485
rect 3764 7451 3798 7485
rect 3832 7451 3866 7485
rect 3900 7451 3934 7485
rect 3968 7451 4002 7485
rect 4036 7451 4070 7485
rect 4104 7451 4138 7485
rect 4172 7451 4206 7485
rect 4240 7451 4274 7485
rect 4308 7451 4342 7485
rect 4376 7451 4410 7485
rect 4444 7451 4478 7485
rect 4512 7451 4546 7485
rect 4580 7451 4614 7485
rect 4648 7451 4682 7485
rect 4716 7451 4750 7485
rect 4784 7451 4818 7485
rect 4852 7451 4886 7485
rect 4920 7451 4954 7485
rect 4988 7451 5022 7485
rect 5056 7451 5090 7485
rect 5124 7451 5158 7485
rect 5192 7451 5226 7485
rect 5260 7451 5294 7485
rect 5328 7451 5362 7485
rect 5396 7451 5430 7485
rect 5464 7451 5498 7485
rect 5532 7451 5566 7485
rect 5600 7451 5634 7485
rect 5668 7451 5702 7485
rect 5736 7451 5770 7485
rect 5804 7451 5838 7485
rect 5872 7451 5906 7485
rect 5940 7451 5974 7485
rect 6008 7451 6042 7485
rect 6076 7451 6110 7485
rect 6144 7451 6178 7485
rect 6212 7451 6246 7485
rect 3508 7329 3542 7363
rect 6316 7329 6350 7363
rect 3508 7261 3542 7295
rect 3508 7193 3542 7227
rect 3508 7125 3542 7159
rect 6316 7261 6350 7295
rect 6316 7193 6350 7227
rect 6316 7125 6350 7159
rect 3508 7057 3542 7091
rect 6316 7057 6350 7091
rect 3508 6989 3542 7023
rect 6316 6989 6350 7023
rect 3508 6921 3542 6955
rect 6316 6921 6350 6955
rect 3508 6853 3542 6887
rect 3508 6785 3542 6819
rect 3508 6717 3542 6751
rect 6316 6853 6350 6887
rect 6316 6785 6350 6819
rect 6316 6717 6350 6751
rect 3508 6649 3542 6683
rect 3508 6581 3542 6615
rect 6316 6649 6350 6683
rect 6316 6581 6350 6615
rect 3508 6513 3542 6547
rect 3508 6445 3542 6479
rect 3508 6377 3542 6411
rect 3508 6309 3542 6343
rect 6316 6445 6350 6479
rect 6316 6377 6350 6411
rect 6316 6309 6350 6343
rect 3508 6241 3542 6275
rect 3508 6173 3542 6207
rect 6316 6241 6350 6275
rect 6316 6173 6350 6207
rect 3508 6105 3542 6139
rect 3508 6037 3542 6071
rect 6316 6105 6350 6139
rect 3508 5969 3542 6003
rect 3508 5901 3542 5935
rect 3508 5833 3542 5867
rect 6316 6037 6350 6071
rect 6316 5969 6350 6003
rect 6316 5901 6350 5935
rect 3508 5765 3542 5799
rect 6316 5833 6350 5867
rect 3508 5697 3542 5731
rect 6316 5765 6350 5799
rect 3508 5629 3542 5663
rect 6316 5697 6350 5731
rect 3508 5561 3542 5595
rect 3508 5493 3542 5527
rect 3508 5425 3542 5459
rect 6316 5629 6350 5663
rect 6316 5561 6350 5595
rect 6316 5493 6350 5527
rect 3508 5357 3542 5391
rect 6316 5425 6350 5459
rect 6316 5357 6350 5391
rect 3508 5289 3542 5323
rect 3508 5221 3542 5255
rect 6316 5289 6350 5323
rect 6316 5221 6350 5255
rect 3508 5153 3542 5187
rect 3508 5085 3542 5119
rect 3508 5017 3542 5051
rect 6316 5153 6350 5187
rect 6316 5085 6350 5119
rect 3508 4949 3542 4983
rect 6316 5017 6350 5051
rect 3508 4881 3542 4915
rect 3508 4813 3542 4847
rect 6316 4881 6350 4915
rect 6316 4813 6350 4847
rect 3508 4745 3542 4779
rect 3508 4677 3542 4711
rect 3508 4609 3542 4643
rect 6316 4745 6350 4779
rect 6316 4677 6350 4711
rect 6316 4609 6350 4643
rect 3508 4541 3542 4575
rect 6316 4541 6350 4575
rect 3508 4473 3542 4507
rect 6316 4473 6350 4507
rect 3508 4405 3542 4439
rect 6316 4405 6350 4439
rect 3508 4337 3542 4371
rect 3508 4269 3542 4303
rect 3508 4201 3542 4235
rect 6316 4337 6350 4371
rect 6316 4269 6350 4303
rect 6316 4201 6350 4235
rect 3508 4133 3542 4167
rect 6316 4133 6350 4167
rect 3628 4011 3662 4045
rect 3696 4011 3730 4045
rect 3764 4011 3798 4045
rect 3832 4011 3866 4045
rect 3900 4011 3934 4045
rect 3968 4011 4002 4045
rect 4036 4011 4070 4045
rect 4104 4011 4138 4045
rect 4172 4011 4206 4045
rect 4240 4011 4274 4045
rect 4308 4011 4342 4045
rect 4376 4011 4410 4045
rect 4444 4011 4478 4045
rect 4512 4011 4546 4045
rect 4580 4011 4614 4045
rect 4648 4011 4682 4045
rect 4716 4011 4750 4045
rect 4784 4011 4818 4045
rect 4852 4011 4886 4045
rect 4920 4011 4954 4045
rect 4988 4011 5022 4045
rect 5056 4011 5090 4045
rect 5124 4011 5158 4045
rect 5192 4011 5226 4045
rect 5260 4011 5294 4045
rect 5328 4011 5362 4045
rect 5396 4011 5430 4045
rect 5464 4011 5498 4045
rect 5532 4011 5566 4045
rect 5600 4011 5634 4045
rect 5668 4011 5702 4045
rect 5736 4011 5770 4045
rect 5804 4011 5838 4045
rect 5872 4011 5906 4045
rect 5940 4011 5974 4045
rect 6008 4011 6042 4045
rect 6076 4011 6110 4045
rect 6144 4011 6178 4045
rect 6212 4011 6246 4045
rect 8364 7040 8398 7074
rect 8432 7040 8466 7074
rect 8500 7040 8534 7074
rect 8568 7040 8602 7074
rect 8636 7040 8670 7074
rect 8704 7040 8738 7074
rect 8772 7040 8806 7074
rect 8840 7040 8874 7074
rect 8908 7040 8942 7074
rect 8976 7040 9010 7074
rect 9044 7040 9078 7074
rect 9112 7040 9146 7074
rect 9180 7040 9214 7074
rect 9248 7040 9282 7074
rect 9316 7040 9350 7074
rect 9384 7040 9418 7074
rect 9452 7040 9486 7074
rect 9520 7040 9554 7074
rect 9588 7040 9622 7074
rect 9656 7040 9690 7074
rect 9724 7040 9758 7074
rect 9792 7040 9826 7074
rect 9860 7040 9894 7074
rect 9928 7040 9962 7074
rect 8244 6918 8278 6952
rect 10020 6918 10054 6952
rect 8244 6850 8278 6884
rect 8244 6782 8278 6816
rect 8244 6714 8278 6748
rect 10020 6850 10054 6884
rect 10020 6782 10054 6816
rect 10020 6714 10054 6748
rect 8244 6646 8278 6680
rect 10020 6646 10054 6680
rect 8244 6578 8278 6612
rect 10020 6578 10054 6612
rect 8244 6510 8278 6544
rect 10020 6510 10054 6544
rect 8244 6442 8278 6476
rect 8244 6374 8278 6408
rect 8244 6306 8278 6340
rect 10020 6442 10054 6476
rect 10020 6374 10054 6408
rect 10020 6306 10054 6340
rect 8244 6238 8278 6272
rect 8244 6170 8278 6204
rect 10020 6238 10054 6272
rect 10020 6170 10054 6204
rect 8244 6102 8278 6136
rect 8244 6034 8278 6068
rect 8244 5966 8278 6000
rect 8244 5898 8278 5932
rect 10020 6034 10054 6068
rect 10020 5966 10054 6000
rect 10020 5898 10054 5932
rect 8244 5830 8278 5864
rect 8244 5762 8278 5796
rect 10020 5830 10054 5864
rect 10020 5762 10054 5796
rect 8244 5694 8278 5728
rect 8244 5626 8278 5660
rect 10020 5694 10054 5728
rect 8244 5558 8278 5592
rect 8244 5490 8278 5524
rect 8244 5422 8278 5456
rect 10020 5626 10054 5660
rect 10020 5558 10054 5592
rect 10020 5490 10054 5524
rect 8244 5354 8278 5388
rect 10020 5422 10054 5456
rect 8244 5286 8278 5320
rect 10020 5354 10054 5388
rect 8244 5218 8278 5252
rect 10020 5286 10054 5320
rect 8244 5150 8278 5184
rect 8244 5082 8278 5116
rect 8244 5014 8278 5048
rect 10020 5218 10054 5252
rect 10020 5150 10054 5184
rect 10020 5082 10054 5116
rect 8244 4946 8278 4980
rect 10020 5014 10054 5048
rect 10020 4946 10054 4980
rect 8244 4878 8278 4912
rect 8244 4810 8278 4844
rect 10020 4878 10054 4912
rect 10020 4810 10054 4844
rect 8244 4742 8278 4776
rect 8244 4674 8278 4708
rect 8244 4606 8278 4640
rect 10020 4742 10054 4776
rect 10020 4674 10054 4708
rect 8244 4538 8278 4572
rect 10020 4606 10054 4640
rect 8244 4470 8278 4504
rect 8244 4402 8278 4436
rect 10020 4470 10054 4504
rect 10020 4402 10054 4436
rect 8244 4334 8278 4368
rect 8244 4266 8278 4300
rect 8244 4198 8278 4232
rect 10020 4334 10054 4368
rect 10020 4266 10054 4300
rect 10020 4198 10054 4232
rect 8244 4130 8278 4164
rect 10020 4130 10054 4164
rect 8364 4018 8398 4052
rect 8432 4018 8466 4052
rect 8500 4018 8534 4052
rect 8568 4018 8602 4052
rect 8636 4018 8670 4052
rect 8704 4018 8738 4052
rect 8772 4018 8806 4052
rect 8840 4018 8874 4052
rect 8908 4018 8942 4052
rect 8976 4018 9010 4052
rect 9044 4018 9078 4052
rect 9112 4018 9146 4052
rect 9180 4018 9214 4052
rect 9248 4018 9282 4052
rect 9316 4018 9350 4052
rect 9384 4018 9418 4052
rect 9452 4018 9486 4052
rect 9520 4018 9554 4052
rect 9588 4018 9622 4052
rect 9656 4018 9690 4052
rect 9724 4018 9758 4052
rect 9792 4018 9826 4052
rect 9860 4018 9894 4052
rect 1518 3956 1552 3990
rect -2202 3814 -2168 3848
rect -2134 3814 -2100 3848
rect -2066 3814 -2032 3848
rect -1998 3814 -1964 3848
rect -1930 3814 -1896 3848
rect -1862 3814 -1828 3848
rect -1794 3814 -1760 3848
rect -1726 3814 -1692 3848
rect -1658 3814 -1624 3848
rect -1590 3814 -1556 3848
rect -1522 3814 -1488 3848
rect -1454 3814 -1420 3848
rect -1386 3814 -1352 3848
rect -1318 3814 -1284 3848
rect -1250 3814 -1216 3848
rect -1182 3814 -1148 3848
rect -1114 3814 -1080 3848
rect -1046 3814 -1012 3848
rect -978 3814 -944 3848
rect -910 3814 -876 3848
rect -842 3814 -808 3848
rect -774 3814 -740 3848
rect -706 3814 -672 3848
rect -638 3814 -604 3848
rect -570 3814 -536 3848
rect -502 3814 -468 3848
rect -434 3814 -400 3848
rect -366 3814 -332 3848
rect -298 3814 -264 3848
rect -230 3814 -196 3848
rect -162 3814 -128 3848
rect -94 3814 -60 3848
rect -26 3814 8 3848
rect 42 3814 76 3848
rect 110 3814 144 3848
rect 178 3814 212 3848
rect 246 3814 280 3848
rect 314 3814 348 3848
rect 382 3814 416 3848
rect 450 3814 484 3848
rect 518 3814 552 3848
rect 586 3814 620 3848
rect 654 3814 688 3848
rect 722 3814 756 3848
rect 790 3814 824 3848
rect 858 3814 892 3848
rect 926 3814 960 3848
rect 994 3814 1028 3848
rect 1062 3814 1096 3848
rect 1130 3814 1164 3848
rect 1198 3814 1232 3848
rect 1266 3814 1300 3848
rect 1334 3814 1368 3848
rect 1402 3814 1436 3848
<< nsubdiffcont >>
rect 7015 10947 7049 10981
rect 7083 10947 7117 10981
rect 7151 10947 7185 10981
rect 7219 10947 7253 10981
rect 7287 10947 7321 10981
rect 7355 10947 7389 10981
rect 7423 10947 7457 10981
rect 7491 10947 7525 10981
rect 7559 10947 7593 10981
rect 7627 10947 7661 10981
rect 7695 10947 7729 10981
rect 7763 10947 7797 10981
rect 7831 10947 7865 10981
rect 7899 10947 7933 10981
rect 7967 10947 8001 10981
rect 8035 10947 8069 10981
rect 8103 10947 8137 10981
rect 8171 10947 8205 10981
rect 8239 10947 8273 10981
rect 8307 10947 8341 10981
rect 8375 10947 8409 10981
rect 8443 10947 8477 10981
rect 8511 10947 8545 10981
rect 8579 10947 8613 10981
rect -1233 10629 -1199 10663
rect -1165 10629 -1131 10663
rect -1097 10629 -1063 10663
rect -1029 10629 -995 10663
rect -961 10629 -927 10663
rect -893 10629 -859 10663
rect -825 10629 -791 10663
rect -757 10629 -723 10663
rect -689 10629 -655 10663
rect -621 10629 -587 10663
rect -553 10629 -519 10663
rect -485 10629 -451 10663
rect -417 10629 -383 10663
rect -349 10629 -315 10663
rect -281 10629 -247 10663
rect -213 10629 -179 10663
rect -145 10629 -111 10663
rect -77 10629 -43 10663
rect -9 10629 25 10663
rect 59 10629 93 10663
rect 127 10629 161 10663
rect 195 10629 229 10663
rect 263 10629 297 10663
rect 331 10629 365 10663
rect -1353 10517 -1319 10551
rect -1353 10449 -1319 10483
rect 423 10517 457 10551
rect -1353 10381 -1319 10415
rect -1353 10313 -1319 10347
rect 423 10449 457 10483
rect 423 10381 457 10415
rect 423 10313 457 10347
rect -1353 10245 -1319 10279
rect -1353 10177 -1319 10211
rect 423 10245 457 10279
rect -1353 10109 -1319 10143
rect 423 10177 457 10211
rect -1353 10041 -1319 10075
rect 423 10109 457 10143
rect -1353 9973 -1319 10007
rect -1353 9905 -1319 9939
rect -1353 9837 -1319 9871
rect 423 10041 457 10075
rect 423 9973 457 10007
rect 423 9905 457 9939
rect -1353 9769 -1319 9803
rect 423 9837 457 9871
rect 423 9769 457 9803
rect -1353 9701 -1319 9735
rect -1353 9633 -1319 9667
rect 423 9701 457 9735
rect 423 9633 457 9667
rect -1353 9565 -1319 9599
rect -1353 9497 -1319 9531
rect -1353 9429 -1319 9463
rect 423 9565 457 9599
rect 423 9497 457 9531
rect 423 9429 457 9463
rect -1353 9361 -1319 9395
rect -1353 9293 -1319 9327
rect 423 9361 457 9395
rect 423 9293 457 9327
rect -1353 9225 -1319 9259
rect -1353 9157 -1319 9191
rect 423 9225 457 9259
rect -1353 9089 -1319 9123
rect -1353 9021 -1319 9055
rect -1353 8953 -1319 8987
rect 423 9157 457 9191
rect 423 9089 457 9123
rect 423 9021 457 9055
rect -1353 8885 -1319 8919
rect 423 8953 457 8987
rect 423 8885 457 8919
rect -1233 8789 -1199 8823
rect -1165 8789 -1131 8823
rect -1097 8789 -1063 8823
rect -1029 8789 -995 8823
rect -961 8789 -927 8823
rect -893 8789 -859 8823
rect -825 8789 -791 8823
rect -757 8789 -723 8823
rect -689 8789 -655 8823
rect -621 8789 -587 8823
rect -553 8789 -519 8823
rect -485 8789 -451 8823
rect -417 8789 -383 8823
rect -349 8789 -315 8823
rect -281 8789 -247 8823
rect -213 8789 -179 8823
rect -145 8789 -111 8823
rect -77 8789 -43 8823
rect -9 8789 25 8823
rect 59 8789 93 8823
rect 127 8789 161 8823
rect 195 8789 229 8823
rect 263 8789 297 8823
rect 331 8789 365 8823
rect 6895 10835 6929 10869
rect 6895 10767 6929 10801
rect 8671 10835 8705 10869
rect 6895 10699 6929 10733
rect 6895 10631 6929 10665
rect 8671 10767 8705 10801
rect 8671 10699 8705 10733
rect 8671 10631 8705 10665
rect 6895 10563 6929 10597
rect 6895 10495 6929 10529
rect 8671 10563 8705 10597
rect 6895 10427 6929 10461
rect 8671 10495 8705 10529
rect 6895 10359 6929 10393
rect 8671 10427 8705 10461
rect 6895 10291 6929 10325
rect 6895 10223 6929 10257
rect 6895 10155 6929 10189
rect 8671 10359 8705 10393
rect 8671 10291 8705 10325
rect 8671 10223 8705 10257
rect 6895 10087 6929 10121
rect 8671 10155 8705 10189
rect 8671 10087 8705 10121
rect 6895 10019 6929 10053
rect 6895 9951 6929 9985
rect 8671 10019 8705 10053
rect 8671 9951 8705 9985
rect 6895 9883 6929 9917
rect 6895 9815 6929 9849
rect 6895 9747 6929 9781
rect 8671 9883 8705 9917
rect 8671 9815 8705 9849
rect 8671 9747 8705 9781
rect 6895 9679 6929 9713
rect 6895 9611 6929 9645
rect 8671 9679 8705 9713
rect 8671 9611 8705 9645
rect 6895 9543 6929 9577
rect 6895 9475 6929 9509
rect 8671 9543 8705 9577
rect 6895 9407 6929 9441
rect 6895 9339 6929 9373
rect 6895 9271 6929 9305
rect 8671 9475 8705 9509
rect 8671 9407 8705 9441
rect 8671 9339 8705 9373
rect 6895 9203 6929 9237
rect 8671 9271 8705 9305
rect 8671 9203 8705 9237
rect 6895 9135 6929 9169
rect 6895 9067 6929 9101
rect 8671 9135 8705 9169
rect 8671 9067 8705 9101
rect 6895 8999 6929 9033
rect 6895 8931 6929 8965
rect 6895 8863 6929 8897
rect 8671 8999 8705 9033
rect 8671 8931 8705 8965
rect 8671 8863 8705 8897
rect 6895 8795 6929 8829
rect 6895 8727 6929 8761
rect 8671 8795 8705 8829
rect 8671 8727 8705 8761
rect 6895 8659 6929 8693
rect 6895 8591 6929 8625
rect 8671 8659 8705 8693
rect 6895 8523 6929 8557
rect 6895 8455 6929 8489
rect 6895 8387 6929 8421
rect 8671 8591 8705 8625
rect 8671 8523 8705 8557
rect 8671 8455 8705 8489
rect 6895 8319 6929 8353
rect 8671 8387 8705 8421
rect 6895 8251 6929 8285
rect 8671 8319 8705 8353
rect 6895 8183 6929 8217
rect 8671 8251 8705 8285
rect 8671 8183 8705 8217
rect 6895 8115 6929 8149
rect 6895 8047 6929 8081
rect 6895 7979 6929 8013
rect 8671 8115 8705 8149
rect 8671 8047 8705 8081
rect 6895 7911 6929 7945
rect 8671 7979 8705 8013
rect 8671 7911 8705 7945
rect 7015 7799 7049 7833
rect 7083 7799 7117 7833
rect 7151 7799 7185 7833
rect 7219 7799 7253 7833
rect 7287 7799 7321 7833
rect 7355 7799 7389 7833
rect 7423 7799 7457 7833
rect 7491 7799 7525 7833
rect 7559 7799 7593 7833
rect 7627 7799 7661 7833
rect 7695 7799 7729 7833
rect 7763 7799 7797 7833
rect 7831 7799 7865 7833
rect 7899 7799 7933 7833
rect 7967 7799 8001 7833
rect 8035 7799 8069 7833
rect 8103 7799 8137 7833
rect 8171 7799 8205 7833
rect 8239 7799 8273 7833
rect 8307 7799 8341 7833
rect 8375 7799 8409 7833
rect 8443 7799 8477 7833
rect 8511 7799 8545 7833
rect 8579 7799 8613 7833
<< poly >>
rect 3129 10771 3329 10787
rect 3129 10737 3178 10771
rect 3212 10737 3246 10771
rect 3280 10737 3329 10771
rect 3129 10699 3329 10737
rect 3387 10771 3587 10787
rect 3387 10737 3436 10771
rect 3470 10737 3504 10771
rect 3538 10737 3587 10771
rect 3387 10699 3587 10737
rect 3645 10771 3845 10787
rect 3645 10737 3694 10771
rect 3728 10737 3762 10771
rect 3796 10737 3845 10771
rect 3645 10699 3845 10737
rect 3903 10699 4103 10787
rect 4161 10699 4361 10787
rect 4419 10771 4619 10787
rect 4419 10737 4468 10771
rect 4502 10737 4536 10771
rect 4570 10737 4619 10771
rect 4419 10699 4619 10737
rect 4677 10771 4877 10787
rect 4677 10737 4726 10771
rect 4760 10737 4794 10771
rect 4828 10737 4877 10771
rect 4677 10699 4877 10737
rect 4935 10771 5135 10787
rect 4935 10737 4984 10771
rect 5018 10737 5052 10771
rect 5086 10737 5135 10771
rect 4935 10699 5135 10737
rect -1193 10561 -993 10577
rect -1193 10527 -1144 10561
rect -1110 10527 -1076 10561
rect -1042 10527 -993 10561
rect -1193 10480 -993 10527
rect -935 10480 -735 10577
rect -677 10480 -477 10577
rect -419 10480 -219 10577
rect -161 10480 39 10577
rect 97 10561 297 10577
rect 97 10527 146 10561
rect 180 10527 214 10561
rect 248 10527 297 10561
rect 97 10480 297 10527
rect -1193 10233 -993 10280
rect -1193 10199 -1144 10233
rect -1110 10199 -1076 10233
rect -1042 10199 -993 10233
rect -1193 10183 -993 10199
rect -935 10233 -735 10280
rect -935 10199 -886 10233
rect -852 10199 -818 10233
rect -784 10199 -735 10233
rect -935 10183 -735 10199
rect -677 10233 -477 10280
rect -677 10199 -628 10233
rect -594 10199 -560 10233
rect -526 10199 -477 10233
rect -677 10183 -477 10199
rect -419 10233 -219 10280
rect -419 10199 -370 10233
rect -336 10199 -302 10233
rect -268 10199 -219 10233
rect -419 10183 -219 10199
rect -161 10233 39 10280
rect -161 10199 -112 10233
rect -78 10199 -44 10233
rect -10 10199 39 10233
rect -161 10183 39 10199
rect 97 10233 297 10280
rect 97 10199 146 10233
rect 180 10199 214 10233
rect 248 10199 297 10233
rect 97 10183 297 10199
rect -1193 10125 -993 10141
rect -1193 10091 -1144 10125
rect -1110 10091 -1076 10125
rect -1042 10091 -993 10125
rect -1193 10044 -993 10091
rect -935 10125 -735 10141
rect -935 10091 -886 10125
rect -852 10091 -818 10125
rect -784 10091 -735 10125
rect -935 10044 -735 10091
rect -677 10125 -477 10141
rect -677 10091 -628 10125
rect -594 10091 -560 10125
rect -526 10091 -477 10125
rect -677 10044 -477 10091
rect -419 10125 -219 10141
rect -419 10091 -370 10125
rect -336 10091 -302 10125
rect -268 10091 -219 10125
rect -419 10044 -219 10091
rect -161 10125 39 10141
rect -161 10091 -112 10125
rect -78 10091 -44 10125
rect -10 10091 39 10125
rect -161 10044 39 10091
rect 97 10125 297 10141
rect 97 10091 146 10125
rect 180 10091 214 10125
rect 248 10091 297 10125
rect 97 10044 297 10091
rect -1193 9797 -993 9844
rect -1193 9763 -1144 9797
rect -1110 9763 -1076 9797
rect -1042 9763 -993 9797
rect -1193 9747 -993 9763
rect -935 9747 -735 9844
rect -677 9747 -477 9844
rect -419 9747 -219 9844
rect -161 9747 39 9844
rect 97 9797 297 9844
rect 97 9763 146 9797
rect 180 9763 214 9797
rect 248 9763 297 9797
rect 97 9747 297 9763
rect -1193 9689 -993 9705
rect -1193 9655 -1144 9689
rect -1110 9655 -1076 9689
rect -1042 9655 -993 9689
rect -1193 9608 -993 9655
rect -935 9608 -735 9705
rect -677 9608 -477 9705
rect -419 9608 -219 9705
rect -161 9608 39 9705
rect 97 9689 297 9705
rect 97 9655 146 9689
rect 180 9655 214 9689
rect 248 9655 297 9689
rect 97 9608 297 9655
rect -1193 9361 -993 9408
rect -1193 9327 -1144 9361
rect -1110 9327 -1076 9361
rect -1042 9327 -993 9361
rect -1193 9311 -993 9327
rect -935 9361 -735 9408
rect -935 9327 -886 9361
rect -852 9327 -818 9361
rect -784 9327 -735 9361
rect -935 9311 -735 9327
rect -677 9361 -477 9408
rect -677 9327 -628 9361
rect -594 9327 -560 9361
rect -526 9327 -477 9361
rect -677 9311 -477 9327
rect -419 9361 -219 9408
rect -419 9327 -370 9361
rect -336 9327 -302 9361
rect -268 9327 -219 9361
rect -419 9311 -219 9327
rect -161 9361 39 9408
rect -161 9327 -112 9361
rect -78 9327 -44 9361
rect -10 9327 39 9361
rect -161 9311 39 9327
rect 97 9361 297 9408
rect 97 9327 146 9361
rect 180 9327 214 9361
rect 248 9327 297 9361
rect 97 9311 297 9327
rect -1193 9253 -993 9269
rect -1193 9219 -1144 9253
rect -1110 9219 -1076 9253
rect -1042 9219 -993 9253
rect -1193 9172 -993 9219
rect -935 9253 -735 9269
rect -935 9219 -886 9253
rect -852 9219 -818 9253
rect -784 9219 -735 9253
rect -935 9172 -735 9219
rect -677 9253 -477 9269
rect -677 9219 -628 9253
rect -594 9219 -560 9253
rect -526 9219 -477 9253
rect -677 9172 -477 9219
rect -419 9253 -219 9269
rect -419 9219 -370 9253
rect -336 9219 -302 9253
rect -268 9219 -219 9253
rect -419 9172 -219 9219
rect -161 9253 39 9269
rect -161 9219 -112 9253
rect -78 9219 -44 9253
rect -10 9219 39 9253
rect -161 9172 39 9219
rect 97 9253 297 9269
rect 97 9219 146 9253
rect 180 9219 214 9253
rect 248 9219 297 9253
rect 97 9172 297 9219
rect -1193 8925 -993 8972
rect -1193 8891 -1144 8925
rect -1110 8891 -1076 8925
rect -1042 8891 -993 8925
rect -1193 8875 -993 8891
rect -935 8875 -735 8972
rect -677 8875 -477 8972
rect -419 8875 -219 8972
rect -161 8875 39 8972
rect 97 8925 297 8972
rect 97 8891 146 8925
rect 180 8891 214 8925
rect 248 8891 297 8925
rect 97 8875 297 8891
rect 3129 10461 3329 10499
rect 3129 10427 3178 10461
rect 3212 10427 3246 10461
rect 3280 10427 3329 10461
rect 3129 10411 3329 10427
rect 3387 10411 3587 10499
rect 3645 10411 3845 10499
rect 3903 10461 4103 10499
rect 3903 10427 3952 10461
rect 3986 10427 4020 10461
rect 4054 10427 4103 10461
rect 3903 10411 4103 10427
rect 4161 10461 4361 10499
rect 4161 10427 4210 10461
rect 4244 10427 4278 10461
rect 4312 10427 4361 10461
rect 4161 10411 4361 10427
rect 4419 10411 4619 10499
rect 4677 10411 4877 10499
rect 4935 10458 5135 10499
rect 4935 10424 4984 10458
rect 5018 10424 5052 10458
rect 5086 10424 5135 10458
rect 4935 10411 5135 10424
rect 3129 10353 3329 10369
rect 3129 10319 3178 10353
rect 3212 10319 3246 10353
rect 3280 10319 3329 10353
rect 3129 10281 3329 10319
rect 3387 10281 3587 10369
rect 3645 10281 3845 10369
rect 3903 10353 4103 10369
rect 3903 10319 3952 10353
rect 3986 10319 4020 10353
rect 4054 10319 4103 10353
rect 3903 10281 4103 10319
rect 4161 10353 4361 10369
rect 4161 10319 4210 10353
rect 4244 10319 4278 10353
rect 4312 10319 4361 10353
rect 4161 10281 4361 10319
rect 4419 10281 4619 10369
rect 4677 10281 4877 10369
rect 4935 10353 5135 10369
rect 4935 10319 4984 10353
rect 5018 10319 5052 10353
rect 5086 10319 5135 10353
rect 4935 10281 5135 10319
rect 3129 10043 3329 10081
rect 3129 10009 3178 10043
rect 3212 10009 3246 10043
rect 3280 10009 3329 10043
rect 3129 9993 3329 10009
rect 3387 10043 3587 10081
rect 3387 10009 3436 10043
rect 3470 10009 3504 10043
rect 3538 10009 3587 10043
rect 3387 9993 3587 10009
rect 3645 10043 3845 10081
rect 3645 10009 3694 10043
rect 3728 10009 3762 10043
rect 3796 10009 3845 10043
rect 3645 9993 3845 10009
rect 3903 9993 4103 10081
rect 4161 9993 4361 10081
rect 4419 10043 4619 10081
rect 4419 10009 4468 10043
rect 4502 10009 4536 10043
rect 4570 10009 4619 10043
rect 4419 9993 4619 10009
rect 4677 10043 4877 10081
rect 4677 10009 4726 10043
rect 4760 10009 4794 10043
rect 4828 10009 4877 10043
rect 4677 9993 4877 10009
rect 4935 10043 5135 10081
rect 4935 10009 4984 10043
rect 5018 10009 5052 10043
rect 5086 10009 5135 10043
rect 4935 9993 5135 10009
rect 3129 9935 3329 9951
rect 3129 9901 3178 9935
rect 3212 9901 3246 9935
rect 3280 9901 3329 9935
rect 3129 9863 3329 9901
rect 3387 9935 3587 9951
rect 3387 9901 3436 9935
rect 3470 9901 3504 9935
rect 3538 9901 3587 9935
rect 3387 9863 3587 9901
rect 3645 9935 3845 9951
rect 3645 9901 3694 9935
rect 3728 9901 3762 9935
rect 3796 9901 3845 9935
rect 3645 9863 3845 9901
rect 3903 9863 4103 9951
rect 4161 9863 4361 9951
rect 4419 9935 4619 9951
rect 4419 9901 4468 9935
rect 4502 9901 4536 9935
rect 4570 9901 4619 9935
rect 4419 9863 4619 9901
rect 4677 9935 4877 9951
rect 4677 9901 4726 9935
rect 4760 9901 4794 9935
rect 4828 9901 4877 9935
rect 4677 9863 4877 9901
rect 4935 9935 5135 9951
rect 4935 9901 4984 9935
rect 5018 9901 5052 9935
rect 5086 9901 5135 9935
rect 4935 9863 5135 9901
rect 3129 9625 3329 9663
rect 3129 9591 3178 9625
rect 3212 9591 3246 9625
rect 3280 9591 3329 9625
rect 3129 9575 3329 9591
rect 3387 9575 3587 9663
rect 3645 9575 3845 9663
rect 3903 9625 4103 9663
rect 3903 9591 3952 9625
rect 3986 9591 4020 9625
rect 4054 9591 4103 9625
rect 3903 9575 4103 9591
rect 4161 9625 4361 9663
rect 4161 9591 4210 9625
rect 4244 9591 4278 9625
rect 4312 9591 4361 9625
rect 4161 9575 4361 9591
rect 4419 9575 4619 9663
rect 4677 9575 4877 9663
rect 4935 9622 5135 9663
rect 4935 9588 4984 9622
rect 5018 9588 5052 9622
rect 5086 9588 5135 9622
rect 4935 9575 5135 9588
rect 3129 9517 3329 9533
rect 3129 9483 3178 9517
rect 3212 9483 3246 9517
rect 3280 9483 3329 9517
rect 3129 9445 3329 9483
rect 3387 9445 3587 9533
rect 3645 9445 3845 9533
rect 3903 9517 4103 9533
rect 3903 9483 3952 9517
rect 3986 9483 4020 9517
rect 4054 9483 4103 9517
rect 3903 9445 4103 9483
rect 4161 9517 4361 9533
rect 4161 9483 4210 9517
rect 4244 9483 4278 9517
rect 4312 9483 4361 9517
rect 4161 9445 4361 9483
rect 4419 9445 4619 9533
rect 4677 9445 4877 9533
rect 4935 9517 5135 9533
rect 4935 9483 4984 9517
rect 5018 9483 5052 9517
rect 5086 9483 5135 9517
rect 4935 9445 5135 9483
rect 3129 9207 3329 9245
rect 3129 9173 3178 9207
rect 3212 9173 3246 9207
rect 3280 9173 3329 9207
rect 3129 9157 3329 9173
rect 3387 9207 3587 9245
rect 3387 9173 3436 9207
rect 3470 9173 3504 9207
rect 3538 9173 3587 9207
rect 3387 9157 3587 9173
rect 3645 9207 3845 9245
rect 3645 9173 3694 9207
rect 3728 9173 3762 9207
rect 3796 9173 3845 9207
rect 3645 9157 3845 9173
rect 3903 9157 4103 9245
rect 4161 9157 4361 9245
rect 4419 9207 4619 9245
rect 4419 9173 4468 9207
rect 4502 9173 4536 9207
rect 4570 9173 4619 9207
rect 4419 9157 4619 9173
rect 4677 9207 4877 9245
rect 4677 9173 4726 9207
rect 4760 9173 4794 9207
rect 4828 9173 4877 9207
rect 4677 9157 4877 9173
rect 4935 9204 5135 9245
rect 4935 9170 4984 9204
rect 5018 9170 5052 9204
rect 5086 9170 5135 9204
rect 4935 9157 5135 9170
rect 3129 9095 3329 9111
rect 3129 9061 3178 9095
rect 3212 9061 3246 9095
rect 3280 9061 3329 9095
rect 3129 9023 3329 9061
rect 3387 9095 3587 9111
rect 3387 9061 3436 9095
rect 3470 9061 3504 9095
rect 3538 9061 3587 9095
rect 3387 9023 3587 9061
rect 3645 9095 3845 9111
rect 3645 9061 3694 9095
rect 3728 9061 3762 9095
rect 3796 9061 3845 9095
rect 3645 9023 3845 9061
rect 3903 9023 4103 9111
rect 4161 9023 4361 9111
rect 4419 9095 4619 9111
rect 4419 9061 4468 9095
rect 4502 9061 4536 9095
rect 4570 9061 4619 9095
rect 4419 9023 4619 9061
rect 4677 9095 4877 9111
rect 4677 9061 4726 9095
rect 4760 9061 4794 9095
rect 4828 9061 4877 9095
rect 4677 9023 4877 9061
rect 4935 9095 5135 9111
rect 4935 9061 4984 9095
rect 5018 9061 5052 9095
rect 5086 9061 5135 9095
rect 4935 9023 5135 9061
rect 3129 8785 3329 8823
rect 3129 8751 3178 8785
rect 3212 8751 3246 8785
rect 3280 8751 3329 8785
rect 3129 8735 3329 8751
rect 3387 8735 3587 8823
rect 3645 8735 3845 8823
rect 3903 8785 4103 8823
rect 3903 8751 3952 8785
rect 3986 8751 4020 8785
rect 4054 8751 4103 8785
rect 3903 8735 4103 8751
rect 4161 8785 4361 8823
rect 4161 8751 4210 8785
rect 4244 8751 4278 8785
rect 4312 8751 4361 8785
rect 4161 8735 4361 8751
rect 4419 8735 4619 8823
rect 4677 8735 4877 8823
rect 4935 8782 5135 8823
rect 4935 8748 4984 8782
rect 5018 8748 5052 8782
rect 5086 8748 5135 8782
rect 4935 8735 5135 8748
rect 3129 8673 3329 8689
rect 3129 8639 3178 8673
rect 3212 8639 3246 8673
rect 3280 8639 3329 8673
rect 3129 8601 3329 8639
rect 3387 8601 3587 8689
rect 3645 8601 3845 8689
rect 3903 8673 4103 8689
rect 3903 8639 3952 8673
rect 3986 8639 4020 8673
rect 4054 8639 4103 8673
rect 3903 8601 4103 8639
rect 4161 8673 4361 8689
rect 4161 8639 4210 8673
rect 4244 8639 4278 8673
rect 4312 8639 4361 8673
rect 4161 8601 4361 8639
rect 4419 8601 4619 8689
rect 4677 8601 4877 8689
rect 4935 8673 5135 8689
rect 4935 8639 4984 8673
rect 5018 8639 5052 8673
rect 5086 8639 5135 8673
rect 4935 8601 5135 8639
rect 3129 8363 3329 8401
rect 3129 8329 3178 8363
rect 3212 8329 3246 8363
rect 3280 8329 3329 8363
rect 3129 8313 3329 8329
rect 3387 8363 3587 8401
rect 3387 8329 3436 8363
rect 3470 8329 3504 8363
rect 3538 8329 3587 8363
rect 3387 8313 3587 8329
rect 3645 8363 3845 8401
rect 3645 8329 3694 8363
rect 3728 8329 3762 8363
rect 3796 8329 3845 8363
rect 3645 8313 3845 8329
rect 3903 8313 4103 8401
rect 4161 8313 4361 8401
rect 4419 8363 4619 8401
rect 4419 8329 4468 8363
rect 4502 8329 4536 8363
rect 4570 8329 4619 8363
rect 4419 8313 4619 8329
rect 4677 8363 4877 8401
rect 4677 8329 4726 8363
rect 4760 8329 4794 8363
rect 4828 8329 4877 8363
rect 4677 8313 4877 8329
rect 4935 8363 5135 8401
rect 4935 8329 4984 8363
rect 5018 8329 5052 8363
rect 5086 8329 5135 8363
rect 4935 8313 5135 8329
rect 7055 10879 7255 10895
rect 7055 10845 7104 10879
rect 7138 10845 7172 10879
rect 7206 10845 7255 10879
rect 7055 10798 7255 10845
rect 7313 10798 7513 10895
rect 7571 10798 7771 10895
rect 7829 10798 8029 10895
rect 8087 10798 8287 10895
rect 8345 10879 8545 10895
rect 8345 10845 8394 10879
rect 8428 10845 8462 10879
rect 8496 10845 8545 10879
rect 8345 10798 8545 10845
rect 7055 10551 7255 10598
rect 7055 10517 7104 10551
rect 7138 10517 7172 10551
rect 7206 10517 7255 10551
rect 7055 10501 7255 10517
rect 7313 10551 7513 10598
rect 7313 10517 7362 10551
rect 7396 10517 7430 10551
rect 7464 10517 7513 10551
rect 7313 10501 7513 10517
rect 7571 10551 7771 10598
rect 7571 10517 7620 10551
rect 7654 10517 7688 10551
rect 7722 10517 7771 10551
rect 7571 10501 7771 10517
rect 7829 10551 8029 10598
rect 7829 10517 7878 10551
rect 7912 10517 7946 10551
rect 7980 10517 8029 10551
rect 7829 10501 8029 10517
rect 8087 10551 8287 10598
rect 8087 10517 8136 10551
rect 8170 10517 8204 10551
rect 8238 10517 8287 10551
rect 8087 10501 8287 10517
rect 8345 10551 8545 10598
rect 8345 10517 8394 10551
rect 8428 10517 8462 10551
rect 8496 10517 8545 10551
rect 8345 10501 8545 10517
rect 7055 10443 7255 10459
rect 7055 10409 7104 10443
rect 7138 10409 7172 10443
rect 7206 10409 7255 10443
rect 7055 10362 7255 10409
rect 7313 10443 7513 10459
rect 7313 10409 7362 10443
rect 7396 10409 7430 10443
rect 7464 10409 7513 10443
rect 7313 10362 7513 10409
rect 7571 10443 7771 10459
rect 7571 10409 7620 10443
rect 7654 10409 7688 10443
rect 7722 10409 7771 10443
rect 7571 10362 7771 10409
rect 7829 10443 8029 10459
rect 7829 10409 7878 10443
rect 7912 10409 7946 10443
rect 7980 10409 8029 10443
rect 7829 10362 8029 10409
rect 8087 10443 8287 10459
rect 8087 10409 8136 10443
rect 8170 10409 8204 10443
rect 8238 10409 8287 10443
rect 8087 10362 8287 10409
rect 8345 10443 8545 10459
rect 8345 10409 8394 10443
rect 8428 10409 8462 10443
rect 8496 10409 8545 10443
rect 8345 10362 8545 10409
rect 7055 10115 7255 10162
rect 7055 10081 7104 10115
rect 7138 10081 7172 10115
rect 7206 10081 7255 10115
rect 7055 10065 7255 10081
rect 7313 10065 7513 10162
rect 7571 10065 7771 10162
rect 7829 10065 8029 10162
rect 8087 10065 8287 10162
rect 8345 10115 8545 10162
rect 8345 10081 8394 10115
rect 8428 10081 8462 10115
rect 8496 10081 8545 10115
rect 8345 10065 8545 10081
rect 7055 10007 7255 10023
rect 7055 9973 7104 10007
rect 7138 9973 7172 10007
rect 7206 9973 7255 10007
rect 7055 9926 7255 9973
rect 7313 9926 7513 10023
rect 7571 9926 7771 10023
rect 7829 9926 8029 10023
rect 8087 9926 8287 10023
rect 8345 10007 8545 10023
rect 8345 9973 8394 10007
rect 8428 9973 8462 10007
rect 8496 9973 8545 10007
rect 8345 9926 8545 9973
rect 7055 9679 7255 9726
rect 7055 9645 7104 9679
rect 7138 9645 7172 9679
rect 7206 9645 7255 9679
rect 7055 9629 7255 9645
rect 7313 9679 7513 9726
rect 7313 9645 7362 9679
rect 7396 9645 7430 9679
rect 7464 9645 7513 9679
rect 7313 9629 7513 9645
rect 7571 9679 7771 9726
rect 7571 9645 7620 9679
rect 7654 9645 7688 9679
rect 7722 9645 7771 9679
rect 7571 9629 7771 9645
rect 7829 9679 8029 9726
rect 7829 9645 7878 9679
rect 7912 9645 7946 9679
rect 7980 9645 8029 9679
rect 7829 9629 8029 9645
rect 8087 9679 8287 9726
rect 8087 9645 8136 9679
rect 8170 9645 8204 9679
rect 8238 9645 8287 9679
rect 8087 9629 8287 9645
rect 8345 9679 8545 9726
rect 8345 9645 8394 9679
rect 8428 9645 8462 9679
rect 8496 9645 8545 9679
rect 8345 9629 8545 9645
rect 7055 9571 7255 9587
rect 7055 9537 7104 9571
rect 7138 9537 7172 9571
rect 7206 9537 7255 9571
rect 7055 9490 7255 9537
rect 7313 9571 7513 9587
rect 7313 9537 7362 9571
rect 7396 9537 7430 9571
rect 7464 9537 7513 9571
rect 7313 9490 7513 9537
rect 7571 9571 7771 9587
rect 7571 9537 7620 9571
rect 7654 9537 7688 9571
rect 7722 9537 7771 9571
rect 7571 9490 7771 9537
rect 7829 9571 8029 9587
rect 7829 9537 7878 9571
rect 7912 9537 7946 9571
rect 7980 9537 8029 9571
rect 7829 9490 8029 9537
rect 8087 9571 8287 9587
rect 8087 9537 8136 9571
rect 8170 9537 8204 9571
rect 8238 9537 8287 9571
rect 8087 9490 8287 9537
rect 8345 9571 8545 9587
rect 8345 9537 8394 9571
rect 8428 9537 8462 9571
rect 8496 9537 8545 9571
rect 8345 9490 8545 9537
rect 7055 9243 7255 9290
rect 7055 9209 7104 9243
rect 7138 9209 7172 9243
rect 7206 9209 7255 9243
rect 7055 9193 7255 9209
rect 7313 9193 7513 9290
rect 7571 9193 7771 9290
rect 7829 9193 8029 9290
rect 8087 9193 8287 9290
rect 8345 9243 8545 9290
rect 8345 9209 8394 9243
rect 8428 9209 8462 9243
rect 8496 9209 8545 9243
rect 8345 9193 8545 9209
rect 7055 9135 7255 9151
rect 7055 9101 7104 9135
rect 7138 9101 7172 9135
rect 7206 9101 7255 9135
rect 7055 9054 7255 9101
rect 7313 9054 7513 9151
rect 7571 9054 7771 9151
rect 7829 9054 8029 9151
rect 8087 9054 8287 9151
rect 8345 9135 8545 9151
rect 8345 9101 8394 9135
rect 8428 9101 8462 9135
rect 8496 9101 8545 9135
rect 8345 9054 8545 9101
rect 7055 8807 7255 8854
rect 7055 8773 7104 8807
rect 7138 8773 7172 8807
rect 7206 8773 7255 8807
rect 7055 8757 7255 8773
rect 7313 8807 7513 8854
rect 7313 8773 7362 8807
rect 7396 8773 7430 8807
rect 7464 8773 7513 8807
rect 7313 8757 7513 8773
rect 7571 8807 7771 8854
rect 7571 8773 7620 8807
rect 7654 8773 7688 8807
rect 7722 8773 7771 8807
rect 7571 8757 7771 8773
rect 7829 8807 8029 8854
rect 7829 8773 7878 8807
rect 7912 8773 7946 8807
rect 7980 8773 8029 8807
rect 7829 8757 8029 8773
rect 8087 8807 8287 8854
rect 8087 8773 8136 8807
rect 8170 8773 8204 8807
rect 8238 8773 8287 8807
rect 8087 8757 8287 8773
rect 8345 8807 8545 8854
rect 8345 8773 8394 8807
rect 8428 8773 8462 8807
rect 8496 8773 8545 8807
rect 8345 8757 8545 8773
rect 7055 8699 7255 8715
rect 7055 8665 7104 8699
rect 7138 8665 7172 8699
rect 7206 8665 7255 8699
rect 7055 8618 7255 8665
rect 7313 8699 7513 8715
rect 7313 8665 7362 8699
rect 7396 8665 7430 8699
rect 7464 8665 7513 8699
rect 7313 8618 7513 8665
rect 7571 8699 7771 8715
rect 7571 8665 7620 8699
rect 7654 8665 7688 8699
rect 7722 8665 7771 8699
rect 7571 8618 7771 8665
rect 7829 8699 8029 8715
rect 7829 8665 7878 8699
rect 7912 8665 7946 8699
rect 7980 8665 8029 8699
rect 7829 8618 8029 8665
rect 8087 8699 8287 8715
rect 8087 8665 8136 8699
rect 8170 8665 8204 8699
rect 8238 8665 8287 8699
rect 8087 8618 8287 8665
rect 8345 8699 8545 8715
rect 8345 8665 8394 8699
rect 8428 8665 8462 8699
rect 8496 8665 8545 8699
rect 8345 8618 8545 8665
rect 7055 8371 7255 8418
rect 7055 8337 7104 8371
rect 7138 8337 7172 8371
rect 7206 8337 7255 8371
rect 7055 8321 7255 8337
rect 7313 8321 7513 8418
rect 7571 8321 7771 8418
rect 7829 8321 8029 8418
rect 8087 8321 8287 8418
rect 8345 8371 8545 8418
rect 8345 8337 8394 8371
rect 8428 8337 8462 8371
rect 8496 8337 8545 8371
rect 8345 8321 8545 8337
rect 7055 8263 7255 8279
rect 7055 8229 7104 8263
rect 7138 8229 7172 8263
rect 7206 8229 7255 8263
rect 7055 8182 7255 8229
rect 7313 8263 7513 8279
rect 7313 8229 7362 8263
rect 7396 8229 7430 8263
rect 7464 8229 7513 8263
rect 7313 8182 7513 8229
rect 7571 8263 7771 8279
rect 7571 8229 7620 8263
rect 7654 8229 7688 8263
rect 7722 8229 7771 8263
rect 7571 8182 7771 8229
rect 7829 8263 8029 8279
rect 7829 8229 7878 8263
rect 7912 8229 7946 8263
rect 7980 8229 8029 8263
rect 7829 8182 8029 8229
rect 8087 8263 8287 8279
rect 8087 8229 8136 8263
rect 8170 8229 8204 8263
rect 8238 8229 8287 8263
rect 8087 8182 8287 8229
rect 8345 8263 8545 8279
rect 8345 8229 8394 8263
rect 8428 8229 8462 8263
rect 8496 8229 8545 8263
rect 8345 8182 8545 8229
rect -2162 8022 -1962 8038
rect -2162 7988 -2113 8022
rect -2079 7988 -2045 8022
rect -2011 7988 -1962 8022
rect -2162 7950 -1962 7988
rect -1904 8022 -1704 8038
rect -1904 7988 -1855 8022
rect -1821 7988 -1787 8022
rect -1753 7988 -1704 8022
rect -1904 7950 -1704 7988
rect -1646 8022 -1446 8038
rect -1646 7988 -1597 8022
rect -1563 7988 -1529 8022
rect -1495 7988 -1446 8022
rect -1646 7950 -1446 7988
rect -1388 8022 -1188 8038
rect -1388 7988 -1339 8022
rect -1305 7988 -1271 8022
rect -1237 7988 -1188 8022
rect -1388 7950 -1188 7988
rect -1130 8022 -930 8038
rect -1130 7988 -1081 8022
rect -1047 7988 -1013 8022
rect -979 7988 -930 8022
rect -1130 7950 -930 7988
rect -872 8022 -672 8038
rect -872 7988 -823 8022
rect -789 7988 -755 8022
rect -721 7988 -672 8022
rect -872 7950 -672 7988
rect -614 8022 -414 8038
rect -614 7988 -565 8022
rect -531 7988 -497 8022
rect -463 7988 -414 8022
rect -614 7950 -414 7988
rect -356 8022 -156 8038
rect -356 7988 -307 8022
rect -273 7988 -239 8022
rect -205 7988 -156 8022
rect -356 7950 -156 7988
rect -98 8022 102 8038
rect -98 7988 -49 8022
rect -15 7988 19 8022
rect 53 7988 102 8022
rect -98 7950 102 7988
rect 160 8022 360 8038
rect 160 7988 209 8022
rect 243 7988 277 8022
rect 311 7988 360 8022
rect 160 7950 360 7988
rect 418 8022 618 8038
rect 418 7988 467 8022
rect 501 7988 535 8022
rect 569 7988 618 8022
rect 418 7950 618 7988
rect 676 8022 876 8038
rect 676 7988 725 8022
rect 759 7988 793 8022
rect 827 7988 876 8022
rect 676 7950 876 7988
rect 934 8022 1134 8038
rect 934 7988 983 8022
rect 1017 7988 1051 8022
rect 1085 7988 1134 8022
rect 934 7950 1134 7988
rect 1192 8022 1392 8038
rect 1192 7988 1241 8022
rect 1275 7988 1309 8022
rect 1343 7988 1392 8022
rect 1192 7950 1392 7988
rect 7055 7935 7255 7982
rect 7055 7901 7104 7935
rect 7138 7901 7172 7935
rect 7206 7901 7255 7935
rect 7055 7885 7255 7901
rect 7313 7885 7513 7982
rect 7571 7885 7771 7982
rect 7829 7885 8029 7982
rect 8087 7885 8287 7982
rect 8345 7935 8545 7982
rect 8345 7901 8394 7935
rect 8428 7901 8462 7935
rect 8496 7901 8545 7935
rect 8345 7885 8545 7901
rect -2162 7712 -1962 7750
rect -2162 7678 -2113 7712
rect -2079 7678 -2045 7712
rect -2011 7678 -1962 7712
rect -2162 7662 -1962 7678
rect -1904 7662 -1704 7750
rect -1646 7662 -1446 7750
rect -1388 7662 -1188 7750
rect -1130 7662 -930 7750
rect -872 7662 -672 7750
rect -614 7662 -414 7750
rect -356 7662 -156 7750
rect -98 7662 102 7750
rect 160 7662 360 7750
rect 418 7662 618 7750
rect 676 7662 876 7750
rect 934 7662 1134 7750
rect 1192 7712 1392 7750
rect 1192 7678 1241 7712
rect 1275 7678 1309 7712
rect 1343 7678 1392 7712
rect 1192 7662 1392 7678
rect -2162 7604 -1962 7620
rect -2162 7570 -2113 7604
rect -2079 7570 -2045 7604
rect -2011 7570 -1962 7604
rect -2162 7532 -1962 7570
rect -1904 7604 -1704 7620
rect -1904 7570 -1855 7604
rect -1821 7570 -1787 7604
rect -1753 7570 -1704 7604
rect -1904 7532 -1704 7570
rect -1646 7604 -1446 7620
rect -1646 7570 -1597 7604
rect -1563 7570 -1529 7604
rect -1495 7570 -1446 7604
rect -1646 7532 -1446 7570
rect -1388 7604 -1188 7620
rect -1388 7570 -1339 7604
rect -1305 7570 -1271 7604
rect -1237 7570 -1188 7604
rect -1388 7532 -1188 7570
rect -1130 7604 -930 7620
rect -1130 7570 -1081 7604
rect -1047 7570 -1013 7604
rect -979 7570 -930 7604
rect -1130 7532 -930 7570
rect -872 7532 -672 7620
rect -614 7532 -414 7620
rect -356 7604 -156 7620
rect -356 7570 -307 7604
rect -273 7570 -239 7604
rect -205 7570 -156 7604
rect -356 7532 -156 7570
rect -98 7604 102 7620
rect -98 7570 -49 7604
rect -15 7570 19 7604
rect 53 7570 102 7604
rect -98 7532 102 7570
rect 160 7532 360 7620
rect 418 7532 618 7620
rect 676 7604 876 7620
rect 676 7570 725 7604
rect 759 7570 793 7604
rect 827 7570 876 7604
rect 676 7532 876 7570
rect 934 7604 1134 7620
rect 934 7570 983 7604
rect 1017 7570 1051 7604
rect 1085 7570 1134 7604
rect 934 7532 1134 7570
rect 1192 7604 1392 7620
rect 1192 7570 1241 7604
rect 1275 7570 1309 7604
rect 1343 7570 1392 7604
rect 1192 7532 1392 7570
rect -2162 7294 -1962 7332
rect -2162 7260 -2113 7294
rect -2079 7260 -2045 7294
rect -2011 7260 -1962 7294
rect -2162 7244 -1962 7260
rect -1904 7244 -1704 7332
rect -1646 7244 -1446 7332
rect -1388 7244 -1188 7332
rect -1130 7244 -930 7332
rect -872 7294 -672 7332
rect -872 7260 -823 7294
rect -789 7260 -755 7294
rect -721 7260 -672 7294
rect -872 7244 -672 7260
rect -614 7294 -414 7332
rect -614 7260 -565 7294
rect -531 7260 -497 7294
rect -463 7260 -414 7294
rect -614 7244 -414 7260
rect -356 7244 -156 7332
rect -98 7244 102 7332
rect 160 7294 360 7332
rect 160 7260 209 7294
rect 243 7260 277 7294
rect 311 7260 360 7294
rect 160 7244 360 7260
rect 418 7294 618 7332
rect 418 7260 467 7294
rect 501 7260 535 7294
rect 569 7260 618 7294
rect 418 7244 618 7260
rect 676 7244 876 7332
rect 934 7244 1134 7332
rect 1192 7294 1392 7332
rect 1192 7260 1241 7294
rect 1275 7260 1309 7294
rect 1343 7260 1392 7294
rect 1192 7244 1392 7260
rect -2162 7186 -1962 7202
rect -2162 7152 -2113 7186
rect -2079 7152 -2045 7186
rect -2011 7152 -1962 7186
rect -2162 7114 -1962 7152
rect -1904 7186 -1704 7202
rect -1904 7152 -1855 7186
rect -1821 7152 -1787 7186
rect -1753 7152 -1704 7186
rect -1904 7114 -1704 7152
rect -1646 7186 -1446 7202
rect -1646 7152 -1597 7186
rect -1563 7152 -1529 7186
rect -1495 7152 -1446 7186
rect -1646 7114 -1446 7152
rect -1388 7114 -1188 7202
rect -1130 7114 -930 7202
rect -872 7186 -672 7202
rect -872 7152 -823 7186
rect -789 7152 -755 7186
rect -721 7152 -672 7186
rect -872 7114 -672 7152
rect -614 7186 -414 7202
rect -614 7152 -565 7186
rect -531 7152 -497 7186
rect -463 7152 -414 7186
rect -614 7114 -414 7152
rect -356 7114 -156 7202
rect -98 7114 102 7202
rect 160 7186 360 7202
rect 160 7152 209 7186
rect 243 7152 277 7186
rect 311 7152 360 7186
rect 160 7114 360 7152
rect 418 7186 618 7202
rect 418 7152 467 7186
rect 501 7152 535 7186
rect 569 7152 618 7186
rect 418 7114 618 7152
rect 676 7114 876 7202
rect 934 7114 1134 7202
rect 1192 7186 1392 7202
rect 1192 7152 1241 7186
rect 1275 7152 1309 7186
rect 1343 7152 1392 7186
rect 1192 7114 1392 7152
rect -2162 6876 -1962 6914
rect -2162 6842 -2113 6876
rect -2079 6842 -2045 6876
rect -2011 6842 -1962 6876
rect -2162 6826 -1962 6842
rect -1904 6826 -1704 6914
rect -1646 6826 -1446 6914
rect -1388 6876 -1188 6914
rect -1388 6842 -1339 6876
rect -1305 6842 -1271 6876
rect -1237 6842 -1188 6876
rect -1388 6826 -1188 6842
rect -1130 6876 -930 6914
rect -1130 6842 -1081 6876
rect -1047 6842 -1013 6876
rect -979 6842 -930 6876
rect -1130 6826 -930 6842
rect -872 6826 -672 6914
rect -614 6826 -414 6914
rect -356 6876 -156 6914
rect -356 6842 -307 6876
rect -273 6842 -239 6876
rect -205 6842 -156 6876
rect -356 6826 -156 6842
rect -98 6876 102 6914
rect -98 6842 -49 6876
rect -15 6842 19 6876
rect 53 6842 102 6876
rect -98 6826 102 6842
rect 160 6826 360 6914
rect 418 6826 618 6914
rect 676 6876 876 6914
rect 676 6842 725 6876
rect 759 6842 793 6876
rect 827 6842 876 6876
rect 676 6826 876 6842
rect 934 6876 1134 6914
rect 934 6842 983 6876
rect 1017 6842 1051 6876
rect 1085 6842 1134 6876
rect 934 6826 1134 6842
rect 1192 6876 1392 6914
rect 1192 6842 1241 6876
rect 1275 6842 1309 6876
rect 1343 6842 1392 6876
rect 1192 6826 1392 6842
rect -2162 6768 -1962 6784
rect -2162 6734 -2113 6768
rect -2079 6734 -2045 6768
rect -2011 6734 -1962 6768
rect -2162 6696 -1962 6734
rect -1904 6696 -1704 6784
rect -1646 6696 -1446 6784
rect -1388 6768 -1188 6784
rect -1388 6734 -1339 6768
rect -1305 6734 -1271 6768
rect -1237 6734 -1188 6768
rect -1388 6696 -1188 6734
rect -1130 6768 -930 6784
rect -1130 6734 -1081 6768
rect -1047 6734 -1013 6768
rect -979 6734 -930 6768
rect -1130 6696 -930 6734
rect -872 6696 -672 6784
rect -614 6696 -414 6784
rect -356 6768 -156 6784
rect -356 6734 -307 6768
rect -273 6734 -239 6768
rect -205 6734 -156 6768
rect -356 6696 -156 6734
rect -98 6768 102 6784
rect -98 6734 -49 6768
rect -15 6734 19 6768
rect 53 6734 102 6768
rect -98 6696 102 6734
rect 160 6696 360 6784
rect 418 6696 618 6784
rect 676 6768 876 6784
rect 676 6734 725 6768
rect 759 6734 793 6768
rect 827 6734 876 6768
rect 676 6696 876 6734
rect 934 6768 1134 6784
rect 934 6734 983 6768
rect 1017 6734 1051 6768
rect 1085 6734 1134 6768
rect 934 6696 1134 6734
rect 1192 6768 1392 6784
rect 1192 6734 1241 6768
rect 1275 6734 1309 6768
rect 1343 6734 1392 6768
rect 1192 6696 1392 6734
rect -2162 6458 -1962 6496
rect -2162 6424 -2113 6458
rect -2079 6424 -2045 6458
rect -2011 6424 -1962 6458
rect -2162 6408 -1962 6424
rect -1904 6458 -1704 6496
rect -1904 6424 -1855 6458
rect -1821 6424 -1787 6458
rect -1753 6424 -1704 6458
rect -1904 6408 -1704 6424
rect -1646 6458 -1446 6496
rect -1646 6424 -1597 6458
rect -1563 6424 -1529 6458
rect -1495 6424 -1446 6458
rect -1646 6408 -1446 6424
rect -1388 6408 -1188 6496
rect -1130 6408 -930 6496
rect -872 6458 -672 6496
rect -872 6424 -823 6458
rect -789 6424 -755 6458
rect -721 6424 -672 6458
rect -872 6408 -672 6424
rect -614 6458 -414 6496
rect -614 6424 -565 6458
rect -531 6424 -497 6458
rect -463 6424 -414 6458
rect -614 6408 -414 6424
rect -356 6408 -156 6496
rect -98 6408 102 6496
rect 160 6458 360 6496
rect 160 6424 209 6458
rect 243 6424 277 6458
rect 311 6424 360 6458
rect 160 6408 360 6424
rect 418 6458 618 6496
rect 418 6424 467 6458
rect 501 6424 535 6458
rect 569 6424 618 6458
rect 418 6408 618 6424
rect 676 6408 876 6496
rect 934 6408 1134 6496
rect 1192 6458 1392 6496
rect 1192 6424 1241 6458
rect 1275 6424 1309 6458
rect 1343 6424 1392 6458
rect 1192 6408 1392 6424
rect -2162 6350 -1962 6366
rect -2162 6316 -2113 6350
rect -2079 6316 -2045 6350
rect -2011 6316 -1962 6350
rect -2162 6278 -1962 6316
rect -1904 6350 -1704 6366
rect -1904 6316 -1855 6350
rect -1821 6316 -1787 6350
rect -1753 6316 -1704 6350
rect -1904 6278 -1704 6316
rect -1646 6350 -1446 6366
rect -1646 6316 -1597 6350
rect -1563 6316 -1529 6350
rect -1495 6316 -1446 6350
rect -1646 6278 -1446 6316
rect -1388 6278 -1188 6366
rect -1130 6278 -930 6366
rect -872 6350 -672 6366
rect -872 6316 -823 6350
rect -789 6316 -755 6350
rect -721 6316 -672 6350
rect -872 6278 -672 6316
rect -614 6350 -414 6366
rect -614 6316 -565 6350
rect -531 6316 -497 6350
rect -463 6316 -414 6350
rect -614 6278 -414 6316
rect -356 6278 -156 6366
rect -98 6278 102 6366
rect 160 6350 360 6366
rect 160 6316 209 6350
rect 243 6316 277 6350
rect 311 6316 360 6350
rect 160 6278 360 6316
rect 418 6350 618 6366
rect 418 6316 467 6350
rect 501 6316 535 6350
rect 569 6316 618 6350
rect 418 6278 618 6316
rect 676 6278 876 6366
rect 934 6278 1134 6366
rect 1192 6350 1392 6366
rect 1192 6316 1241 6350
rect 1275 6316 1309 6350
rect 1343 6316 1392 6350
rect 1192 6278 1392 6316
rect -2162 6040 -1962 6078
rect -2162 6006 -2113 6040
rect -2079 6006 -2045 6040
rect -2011 6006 -1962 6040
rect -2162 5990 -1962 6006
rect -1904 5990 -1704 6078
rect -1646 5990 -1446 6078
rect -1388 6040 -1188 6078
rect -1388 6006 -1339 6040
rect -1305 6006 -1271 6040
rect -1237 6006 -1188 6040
rect -1388 5990 -1188 6006
rect -1130 6040 -930 6078
rect -1130 6006 -1081 6040
rect -1047 6006 -1013 6040
rect -979 6006 -930 6040
rect -1130 5990 -930 6006
rect -872 5990 -672 6078
rect -614 5990 -414 6078
rect -356 6040 -156 6078
rect -356 6006 -307 6040
rect -273 6006 -239 6040
rect -205 6006 -156 6040
rect -356 5990 -156 6006
rect -98 6040 102 6078
rect -98 6006 -49 6040
rect -15 6006 19 6040
rect 53 6006 102 6040
rect -98 5990 102 6006
rect 160 5990 360 6078
rect 418 5990 618 6078
rect 676 6040 876 6078
rect 676 6006 725 6040
rect 759 6006 793 6040
rect 827 6006 876 6040
rect 676 5990 876 6006
rect 934 6040 1134 6078
rect 934 6006 983 6040
rect 1017 6006 1051 6040
rect 1085 6006 1134 6040
rect 934 5990 1134 6006
rect 1192 6040 1392 6078
rect 1192 6006 1241 6040
rect 1275 6006 1309 6040
rect 1343 6006 1392 6040
rect 1192 5990 1392 6006
rect -2162 5932 -1962 5948
rect -2162 5898 -2113 5932
rect -2079 5898 -2045 5932
rect -2011 5898 -1962 5932
rect -2162 5860 -1962 5898
rect -1904 5860 -1704 5948
rect -1646 5860 -1446 5948
rect -1388 5932 -1188 5948
rect -1388 5898 -1339 5932
rect -1305 5898 -1271 5932
rect -1237 5898 -1188 5932
rect -1388 5860 -1188 5898
rect -1130 5932 -930 5948
rect -1130 5898 -1081 5932
rect -1047 5898 -1013 5932
rect -979 5898 -930 5932
rect -1130 5860 -930 5898
rect -872 5860 -672 5948
rect -614 5860 -414 5948
rect -356 5932 -156 5948
rect -356 5898 -307 5932
rect -273 5898 -239 5932
rect -205 5898 -156 5932
rect -356 5860 -156 5898
rect -98 5932 102 5948
rect -98 5898 -49 5932
rect -15 5898 19 5932
rect 53 5898 102 5932
rect -98 5860 102 5898
rect 160 5860 360 5948
rect 418 5860 618 5948
rect 676 5932 876 5948
rect 676 5898 725 5932
rect 759 5898 793 5932
rect 827 5898 876 5932
rect 676 5860 876 5898
rect 934 5932 1134 5948
rect 934 5898 983 5932
rect 1017 5898 1051 5932
rect 1085 5898 1134 5932
rect 934 5860 1134 5898
rect 1192 5932 1392 5948
rect 1192 5898 1241 5932
rect 1275 5898 1309 5932
rect 1343 5898 1392 5932
rect 1192 5860 1392 5898
rect -2162 5622 -1962 5660
rect -2162 5588 -2113 5622
rect -2079 5588 -2045 5622
rect -2011 5588 -1962 5622
rect -2162 5572 -1962 5588
rect -1904 5622 -1704 5660
rect -1904 5588 -1855 5622
rect -1821 5588 -1787 5622
rect -1753 5588 -1704 5622
rect -1904 5572 -1704 5588
rect -1646 5622 -1446 5660
rect -1646 5588 -1597 5622
rect -1563 5588 -1529 5622
rect -1495 5588 -1446 5622
rect -1646 5572 -1446 5588
rect -1388 5572 -1188 5660
rect -1130 5572 -930 5660
rect -872 5622 -672 5660
rect -872 5588 -823 5622
rect -789 5588 -755 5622
rect -721 5588 -672 5622
rect -872 5572 -672 5588
rect -614 5622 -414 5660
rect -614 5588 -565 5622
rect -531 5588 -497 5622
rect -463 5588 -414 5622
rect -614 5572 -414 5588
rect -356 5572 -156 5660
rect -98 5572 102 5660
rect 160 5622 360 5660
rect 160 5588 209 5622
rect 243 5588 277 5622
rect 311 5588 360 5622
rect 160 5572 360 5588
rect 418 5622 618 5660
rect 418 5588 467 5622
rect 501 5588 535 5622
rect 569 5588 618 5622
rect 418 5572 618 5588
rect 676 5572 876 5660
rect 934 5572 1134 5660
rect 1192 5622 1392 5660
rect 1192 5588 1241 5622
rect 1275 5588 1309 5622
rect 1343 5588 1392 5622
rect 1192 5572 1392 5588
rect -2162 5514 -1962 5530
rect -2162 5480 -2113 5514
rect -2079 5480 -2045 5514
rect -2011 5480 -1962 5514
rect -2162 5442 -1962 5480
rect -1904 5514 -1704 5530
rect -1904 5480 -1855 5514
rect -1821 5480 -1787 5514
rect -1753 5480 -1704 5514
rect -1904 5442 -1704 5480
rect -1646 5514 -1446 5530
rect -1646 5480 -1597 5514
rect -1563 5480 -1529 5514
rect -1495 5480 -1446 5514
rect -1646 5442 -1446 5480
rect -1388 5442 -1188 5530
rect -1130 5442 -930 5530
rect -872 5514 -672 5530
rect -872 5480 -823 5514
rect -789 5480 -755 5514
rect -721 5480 -672 5514
rect -872 5442 -672 5480
rect -614 5514 -414 5530
rect -614 5480 -565 5514
rect -531 5480 -497 5514
rect -463 5480 -414 5514
rect -614 5442 -414 5480
rect -356 5442 -156 5530
rect -98 5442 102 5530
rect 160 5514 360 5530
rect 160 5480 209 5514
rect 243 5480 277 5514
rect 311 5480 360 5514
rect 160 5442 360 5480
rect 418 5514 618 5530
rect 418 5480 467 5514
rect 501 5480 535 5514
rect 569 5480 618 5514
rect 418 5442 618 5480
rect 676 5442 876 5530
rect 934 5442 1134 5530
rect 1192 5514 1392 5530
rect 1192 5480 1241 5514
rect 1275 5480 1309 5514
rect 1343 5480 1392 5514
rect 1192 5442 1392 5480
rect -2162 5204 -1962 5242
rect -2162 5170 -2113 5204
rect -2079 5170 -2045 5204
rect -2011 5170 -1962 5204
rect -2162 5154 -1962 5170
rect -1904 5154 -1704 5242
rect -1646 5154 -1446 5242
rect -1388 5204 -1188 5242
rect -1388 5170 -1339 5204
rect -1305 5170 -1271 5204
rect -1237 5170 -1188 5204
rect -1388 5154 -1188 5170
rect -1130 5204 -930 5242
rect -1130 5170 -1081 5204
rect -1047 5170 -1013 5204
rect -979 5170 -930 5204
rect -1130 5154 -930 5170
rect -872 5154 -672 5242
rect -614 5154 -414 5242
rect -356 5204 -156 5242
rect -356 5170 -307 5204
rect -273 5170 -239 5204
rect -205 5170 -156 5204
rect -356 5154 -156 5170
rect -98 5204 102 5242
rect -98 5170 -49 5204
rect -15 5170 19 5204
rect 53 5170 102 5204
rect -98 5154 102 5170
rect 160 5154 360 5242
rect 418 5154 618 5242
rect 676 5204 876 5242
rect 676 5170 725 5204
rect 759 5170 793 5204
rect 827 5170 876 5204
rect 676 5154 876 5170
rect 934 5204 1134 5242
rect 934 5170 983 5204
rect 1017 5170 1051 5204
rect 1085 5170 1134 5204
rect 934 5154 1134 5170
rect 1192 5204 1392 5242
rect 1192 5170 1241 5204
rect 1275 5170 1309 5204
rect 1343 5170 1392 5204
rect 1192 5154 1392 5170
rect -2162 5096 -1962 5112
rect -2162 5062 -2113 5096
rect -2079 5062 -2045 5096
rect -2011 5062 -1962 5096
rect -2162 5024 -1962 5062
rect -1904 5024 -1704 5112
rect -1646 5024 -1446 5112
rect -1388 5096 -1188 5112
rect -1388 5062 -1339 5096
rect -1305 5062 -1271 5096
rect -1237 5062 -1188 5096
rect -1388 5024 -1188 5062
rect -1130 5096 -930 5112
rect -1130 5062 -1081 5096
rect -1047 5062 -1013 5096
rect -979 5062 -930 5096
rect -1130 5024 -930 5062
rect -872 5024 -672 5112
rect -614 5024 -414 5112
rect -356 5096 -156 5112
rect -356 5062 -307 5096
rect -273 5062 -239 5096
rect -205 5062 -156 5096
rect -356 5024 -156 5062
rect -98 5096 102 5112
rect -98 5062 -49 5096
rect -15 5062 19 5096
rect 53 5062 102 5096
rect -98 5024 102 5062
rect 160 5024 360 5112
rect 418 5024 618 5112
rect 676 5096 876 5112
rect 676 5062 725 5096
rect 759 5062 793 5096
rect 827 5062 876 5096
rect 676 5024 876 5062
rect 934 5096 1134 5112
rect 934 5062 983 5096
rect 1017 5062 1051 5096
rect 1085 5062 1134 5096
rect 934 5024 1134 5062
rect 1192 5096 1392 5112
rect 1192 5062 1241 5096
rect 1275 5062 1309 5096
rect 1343 5062 1392 5096
rect 1192 5024 1392 5062
rect -2162 4786 -1962 4824
rect -2162 4752 -2113 4786
rect -2079 4752 -2045 4786
rect -2011 4752 -1962 4786
rect -2162 4736 -1962 4752
rect -1904 4786 -1704 4824
rect -1904 4752 -1855 4786
rect -1821 4752 -1787 4786
rect -1753 4752 -1704 4786
rect -1904 4736 -1704 4752
rect -1646 4786 -1446 4824
rect -1646 4752 -1597 4786
rect -1563 4752 -1529 4786
rect -1495 4752 -1446 4786
rect -1646 4736 -1446 4752
rect -1388 4736 -1188 4824
rect -1130 4736 -930 4824
rect -872 4786 -672 4824
rect -872 4752 -823 4786
rect -789 4752 -755 4786
rect -721 4752 -672 4786
rect -872 4736 -672 4752
rect -614 4786 -414 4824
rect -614 4752 -565 4786
rect -531 4752 -497 4786
rect -463 4752 -414 4786
rect -614 4736 -414 4752
rect -356 4736 -156 4824
rect -98 4736 102 4824
rect 160 4786 360 4824
rect 160 4752 209 4786
rect 243 4752 277 4786
rect 311 4752 360 4786
rect 160 4736 360 4752
rect 418 4786 618 4824
rect 418 4752 467 4786
rect 501 4752 535 4786
rect 569 4752 618 4786
rect 418 4736 618 4752
rect 676 4736 876 4824
rect 934 4736 1134 4824
rect 1192 4786 1392 4824
rect 1192 4752 1241 4786
rect 1275 4752 1309 4786
rect 1343 4752 1392 4786
rect 1192 4736 1392 4752
rect -2162 4678 -1962 4694
rect -2162 4644 -2113 4678
rect -2079 4644 -2045 4678
rect -2011 4644 -1962 4678
rect -2162 4606 -1962 4644
rect -1904 4678 -1704 4694
rect -1904 4644 -1855 4678
rect -1821 4644 -1787 4678
rect -1753 4644 -1704 4678
rect -1904 4606 -1704 4644
rect -1646 4678 -1446 4694
rect -1646 4644 -1597 4678
rect -1563 4644 -1529 4678
rect -1495 4644 -1446 4678
rect -1646 4606 -1446 4644
rect -1388 4606 -1188 4694
rect -1130 4606 -930 4694
rect -872 4678 -672 4694
rect -872 4644 -823 4678
rect -789 4644 -755 4678
rect -721 4644 -672 4678
rect -872 4606 -672 4644
rect -614 4678 -414 4694
rect -614 4644 -565 4678
rect -531 4644 -497 4678
rect -463 4644 -414 4678
rect -614 4606 -414 4644
rect -356 4606 -156 4694
rect -98 4606 102 4694
rect 160 4678 360 4694
rect 160 4644 209 4678
rect 243 4644 277 4678
rect 311 4644 360 4678
rect 160 4606 360 4644
rect 418 4678 618 4694
rect 418 4644 467 4678
rect 501 4644 535 4678
rect 569 4644 618 4678
rect 418 4606 618 4644
rect 676 4678 876 4694
rect 676 4644 725 4678
rect 759 4644 793 4678
rect 827 4644 876 4678
rect 676 4606 876 4644
rect 934 4678 1134 4694
rect 934 4644 983 4678
rect 1017 4644 1051 4678
rect 1085 4644 1134 4678
rect 934 4606 1134 4644
rect 1192 4678 1392 4694
rect 1192 4644 1241 4678
rect 1275 4644 1309 4678
rect 1343 4644 1392 4678
rect 1192 4606 1392 4644
rect -2162 4368 -1962 4406
rect -2162 4334 -2113 4368
rect -2079 4334 -2045 4368
rect -2011 4334 -1962 4368
rect -2162 4318 -1962 4334
rect -1904 4318 -1704 4406
rect -1646 4318 -1446 4406
rect -1388 4368 -1188 4406
rect -1388 4334 -1339 4368
rect -1305 4334 -1271 4368
rect -1237 4334 -1188 4368
rect -1388 4318 -1188 4334
rect -1130 4368 -930 4406
rect -1130 4334 -1081 4368
rect -1047 4334 -1013 4368
rect -979 4334 -930 4368
rect -1130 4318 -930 4334
rect -872 4318 -672 4406
rect -614 4318 -414 4406
rect -356 4368 -156 4406
rect -356 4334 -307 4368
rect -273 4334 -239 4368
rect -205 4334 -156 4368
rect -356 4318 -156 4334
rect -98 4368 102 4406
rect -98 4334 -49 4368
rect -15 4334 19 4368
rect 53 4334 102 4368
rect -98 4318 102 4334
rect 160 4318 360 4406
rect 418 4318 618 4406
rect 676 4318 876 4406
rect 934 4318 1134 4406
rect 1192 4368 1392 4406
rect 1192 4334 1241 4368
rect 1275 4334 1309 4368
rect 1343 4334 1392 4368
rect 1192 4318 1392 4334
rect -2162 4260 -1962 4276
rect -2162 4226 -2113 4260
rect -2079 4226 -2045 4260
rect -2011 4226 -1962 4260
rect -2162 4188 -1962 4226
rect -1904 4260 -1704 4276
rect -1904 4226 -1855 4260
rect -1821 4226 -1787 4260
rect -1753 4226 -1704 4260
rect -1904 4188 -1704 4226
rect -1646 4260 -1446 4276
rect -1646 4226 -1597 4260
rect -1563 4226 -1529 4260
rect -1495 4226 -1446 4260
rect -1646 4188 -1446 4226
rect -1388 4260 -1188 4276
rect -1388 4226 -1339 4260
rect -1305 4226 -1271 4260
rect -1237 4226 -1188 4260
rect -1388 4188 -1188 4226
rect -1130 4260 -930 4276
rect -1130 4226 -1081 4260
rect -1047 4226 -1013 4260
rect -979 4226 -930 4260
rect -1130 4188 -930 4226
rect -872 4260 -672 4276
rect -872 4226 -823 4260
rect -789 4226 -755 4260
rect -721 4226 -672 4260
rect -872 4188 -672 4226
rect -614 4260 -414 4276
rect -614 4226 -565 4260
rect -531 4226 -497 4260
rect -463 4226 -414 4260
rect -614 4188 -414 4226
rect -356 4260 -156 4276
rect -356 4226 -307 4260
rect -273 4226 -239 4260
rect -205 4226 -156 4260
rect -356 4188 -156 4226
rect -98 4260 102 4276
rect -98 4226 -49 4260
rect -15 4226 19 4260
rect 53 4226 102 4260
rect -98 4188 102 4226
rect 160 4260 360 4276
rect 160 4226 209 4260
rect 243 4226 277 4260
rect 311 4226 360 4260
rect 160 4188 360 4226
rect 418 4260 618 4276
rect 418 4226 467 4260
rect 501 4226 535 4260
rect 569 4226 618 4260
rect 418 4188 618 4226
rect 676 4260 876 4276
rect 676 4226 725 4260
rect 759 4226 793 4260
rect 827 4226 876 4260
rect 676 4188 876 4226
rect 934 4260 1134 4276
rect 934 4226 983 4260
rect 1017 4226 1051 4260
rect 1085 4226 1134 4260
rect 934 4188 1134 4226
rect 1192 4260 1392 4276
rect 1192 4226 1241 4260
rect 1275 4226 1309 4260
rect 1343 4226 1392 4260
rect 1192 4188 1392 4226
rect 3668 7383 3868 7399
rect 3668 7349 3717 7383
rect 3751 7349 3785 7383
rect 3819 7349 3868 7383
rect 3668 7311 3868 7349
rect 3926 7383 4126 7399
rect 3926 7349 3975 7383
rect 4009 7349 4043 7383
rect 4077 7349 4126 7383
rect 3926 7311 4126 7349
rect 4184 7383 4384 7399
rect 4184 7349 4233 7383
rect 4267 7349 4301 7383
rect 4335 7349 4384 7383
rect 4184 7311 4384 7349
rect 4442 7383 4642 7399
rect 4442 7349 4491 7383
rect 4525 7349 4559 7383
rect 4593 7349 4642 7383
rect 4442 7311 4642 7349
rect 4700 7383 4900 7399
rect 4700 7349 4749 7383
rect 4783 7349 4817 7383
rect 4851 7349 4900 7383
rect 4700 7311 4900 7349
rect 4958 7383 5158 7399
rect 4958 7349 5007 7383
rect 5041 7349 5075 7383
rect 5109 7349 5158 7383
rect 4958 7311 5158 7349
rect 5216 7383 5416 7399
rect 5216 7349 5265 7383
rect 5299 7349 5333 7383
rect 5367 7349 5416 7383
rect 5216 7311 5416 7349
rect 5474 7383 5674 7399
rect 5474 7349 5523 7383
rect 5557 7349 5591 7383
rect 5625 7349 5674 7383
rect 5474 7311 5674 7349
rect 5732 7383 5932 7399
rect 5732 7349 5781 7383
rect 5815 7349 5849 7383
rect 5883 7349 5932 7383
rect 5732 7311 5932 7349
rect 5990 7383 6190 7399
rect 5990 7349 6039 7383
rect 6073 7349 6107 7383
rect 6141 7349 6190 7383
rect 5990 7311 6190 7349
rect 3668 7073 3868 7111
rect 3668 7039 3717 7073
rect 3751 7039 3785 7073
rect 3819 7039 3868 7073
rect 3668 7023 3868 7039
rect 3926 7023 4126 7111
rect 4184 7023 4384 7111
rect 4442 7023 4642 7111
rect 4700 7023 4900 7111
rect 4958 7023 5158 7111
rect 5216 7023 5416 7111
rect 5474 7023 5674 7111
rect 5732 7023 5932 7111
rect 5990 7073 6190 7111
rect 5990 7039 6039 7073
rect 6073 7039 6107 7073
rect 6141 7039 6190 7073
rect 5990 7023 6190 7039
rect 3668 6965 3868 6981
rect 3668 6931 3717 6965
rect 3751 6931 3785 6965
rect 3819 6931 3868 6965
rect 3668 6893 3868 6931
rect 3926 6965 4126 6981
rect 3926 6931 3975 6965
rect 4009 6931 4043 6965
rect 4077 6931 4126 6965
rect 3926 6893 4126 6931
rect 4184 6965 4384 6981
rect 4184 6931 4233 6965
rect 4267 6931 4301 6965
rect 4335 6931 4384 6965
rect 4184 6893 4384 6931
rect 4442 6893 4642 6981
rect 4700 6893 4900 6981
rect 4958 6965 5158 6981
rect 4958 6931 5007 6965
rect 5041 6931 5075 6965
rect 5109 6931 5158 6965
rect 4958 6893 5158 6931
rect 5216 6965 5416 6981
rect 5216 6931 5265 6965
rect 5299 6931 5333 6965
rect 5367 6931 5416 6965
rect 5216 6893 5416 6931
rect 5474 6893 5674 6981
rect 5732 6893 5932 6981
rect 5990 6965 6190 6981
rect 5990 6931 6039 6965
rect 6073 6931 6107 6965
rect 6141 6931 6190 6965
rect 5990 6893 6190 6931
rect 3668 6655 3868 6693
rect 3668 6621 3717 6655
rect 3751 6621 3785 6655
rect 3819 6621 3868 6655
rect 3668 6605 3868 6621
rect 3926 6605 4126 6693
rect 4184 6605 4384 6693
rect 4442 6655 4642 6693
rect 4442 6621 4491 6655
rect 4525 6621 4559 6655
rect 4593 6621 4642 6655
rect 4442 6605 4642 6621
rect 4700 6655 4900 6693
rect 4700 6621 4749 6655
rect 4783 6621 4817 6655
rect 4851 6621 4900 6655
rect 4700 6605 4900 6621
rect 4958 6605 5158 6693
rect 5216 6605 5416 6693
rect 5474 6655 5674 6693
rect 5474 6621 5523 6655
rect 5557 6621 5591 6655
rect 5625 6621 5674 6655
rect 5474 6605 5674 6621
rect 5732 6655 5932 6693
rect 5732 6621 5781 6655
rect 5815 6621 5849 6655
rect 5883 6621 5932 6655
rect 5732 6605 5932 6621
rect 5990 6655 6190 6693
rect 5990 6621 6039 6655
rect 6073 6621 6107 6655
rect 6141 6621 6190 6655
rect 5990 6605 6190 6621
rect 3668 6547 3868 6563
rect 3668 6513 3717 6547
rect 3751 6513 3785 6547
rect 3819 6513 3868 6547
rect 3668 6475 3868 6513
rect 3926 6475 4126 6563
rect 4184 6475 4384 6563
rect 4442 6547 4642 6563
rect 4442 6513 4491 6547
rect 4525 6513 4559 6547
rect 4593 6513 4642 6547
rect 4442 6475 4642 6513
rect 4700 6547 4900 6563
rect 4700 6513 4749 6547
rect 4783 6513 4817 6547
rect 4851 6513 4900 6547
rect 4700 6475 4900 6513
rect 4958 6475 5158 6563
rect 5216 6475 5416 6563
rect 5474 6547 5674 6563
rect 5474 6513 5523 6547
rect 5557 6513 5591 6547
rect 5625 6513 5674 6547
rect 5474 6475 5674 6513
rect 5732 6547 5932 6563
rect 5732 6513 5781 6547
rect 5815 6513 5849 6547
rect 5883 6513 5932 6547
rect 5732 6475 5932 6513
rect 5990 6547 6190 6563
rect 5990 6513 6039 6547
rect 6073 6513 6107 6547
rect 6141 6513 6190 6547
rect 5990 6475 6190 6513
rect 3668 6237 3868 6275
rect 3668 6203 3717 6237
rect 3751 6203 3785 6237
rect 3819 6203 3868 6237
rect 3668 6187 3868 6203
rect 3926 6237 4126 6275
rect 3926 6203 3975 6237
rect 4009 6203 4043 6237
rect 4077 6203 4126 6237
rect 3926 6187 4126 6203
rect 4184 6237 4384 6275
rect 4184 6203 4233 6237
rect 4267 6203 4301 6237
rect 4335 6203 4384 6237
rect 4184 6187 4384 6203
rect 4442 6187 4642 6275
rect 4700 6187 4900 6275
rect 4958 6237 5158 6275
rect 4958 6203 5007 6237
rect 5041 6203 5075 6237
rect 5109 6203 5158 6237
rect 4958 6187 5158 6203
rect 5216 6237 5416 6275
rect 5216 6203 5265 6237
rect 5299 6203 5333 6237
rect 5367 6203 5416 6237
rect 5216 6187 5416 6203
rect 5474 6187 5674 6275
rect 5732 6187 5932 6275
rect 5990 6237 6190 6275
rect 5990 6203 6039 6237
rect 6073 6203 6107 6237
rect 6141 6203 6190 6237
rect 5990 6187 6190 6203
rect 3668 6129 3868 6145
rect 3668 6095 3717 6129
rect 3751 6095 3785 6129
rect 3819 6095 3868 6129
rect 3668 6057 3868 6095
rect 3926 6129 4126 6145
rect 3926 6095 3975 6129
rect 4009 6095 4043 6129
rect 4077 6095 4126 6129
rect 3926 6057 4126 6095
rect 4184 6129 4384 6145
rect 4184 6095 4233 6129
rect 4267 6095 4301 6129
rect 4335 6095 4384 6129
rect 4184 6057 4384 6095
rect 4442 6057 4642 6145
rect 4700 6057 4900 6145
rect 4958 6129 5158 6145
rect 4958 6095 5007 6129
rect 5041 6095 5075 6129
rect 5109 6095 5158 6129
rect 4958 6057 5158 6095
rect 5216 6129 5416 6145
rect 5216 6095 5265 6129
rect 5299 6095 5333 6129
rect 5367 6095 5416 6129
rect 5216 6057 5416 6095
rect 5474 6057 5674 6145
rect 5732 6057 5932 6145
rect 5990 6129 6190 6145
rect 5990 6095 6039 6129
rect 6073 6095 6107 6129
rect 6141 6095 6190 6129
rect 5990 6057 6190 6095
rect 3668 5819 3868 5857
rect 3668 5785 3717 5819
rect 3751 5785 3785 5819
rect 3819 5785 3868 5819
rect 3668 5769 3868 5785
rect 3926 5769 4126 5857
rect 4184 5769 4384 5857
rect 4442 5819 4642 5857
rect 4442 5785 4491 5819
rect 4525 5785 4559 5819
rect 4593 5785 4642 5819
rect 4442 5769 4642 5785
rect 4700 5819 4900 5857
rect 4700 5785 4749 5819
rect 4783 5785 4817 5819
rect 4851 5785 4900 5819
rect 4700 5769 4900 5785
rect 4958 5769 5158 5857
rect 5216 5769 5416 5857
rect 5474 5819 5674 5857
rect 5474 5785 5523 5819
rect 5557 5785 5591 5819
rect 5625 5785 5674 5819
rect 5474 5769 5674 5785
rect 5732 5819 5932 5857
rect 5732 5785 5781 5819
rect 5815 5785 5849 5819
rect 5883 5785 5932 5819
rect 5732 5769 5932 5785
rect 5990 5819 6190 5857
rect 5990 5785 6039 5819
rect 6073 5785 6107 5819
rect 6141 5785 6190 5819
rect 5990 5769 6190 5785
rect 3668 5711 3868 5727
rect 3668 5677 3717 5711
rect 3751 5677 3785 5711
rect 3819 5677 3868 5711
rect 3668 5639 3868 5677
rect 3926 5639 4126 5727
rect 4184 5639 4384 5727
rect 4442 5711 4642 5727
rect 4442 5677 4491 5711
rect 4525 5677 4559 5711
rect 4593 5677 4642 5711
rect 4442 5639 4642 5677
rect 4700 5711 4900 5727
rect 4700 5677 4749 5711
rect 4783 5677 4817 5711
rect 4851 5677 4900 5711
rect 4700 5639 4900 5677
rect 4958 5639 5158 5727
rect 5216 5639 5416 5727
rect 5474 5711 5674 5727
rect 5474 5677 5523 5711
rect 5557 5677 5591 5711
rect 5625 5677 5674 5711
rect 5474 5639 5674 5677
rect 5732 5711 5932 5727
rect 5732 5677 5781 5711
rect 5815 5677 5849 5711
rect 5883 5677 5932 5711
rect 5732 5639 5932 5677
rect 5990 5711 6190 5727
rect 5990 5677 6039 5711
rect 6073 5677 6107 5711
rect 6141 5677 6190 5711
rect 5990 5639 6190 5677
rect 3668 5401 3868 5439
rect 3668 5367 3717 5401
rect 3751 5367 3785 5401
rect 3819 5367 3868 5401
rect 3668 5351 3868 5367
rect 3926 5401 4126 5439
rect 3926 5367 3975 5401
rect 4009 5367 4043 5401
rect 4077 5367 4126 5401
rect 3926 5351 4126 5367
rect 4184 5401 4384 5439
rect 4184 5367 4233 5401
rect 4267 5367 4301 5401
rect 4335 5367 4384 5401
rect 4184 5351 4384 5367
rect 4442 5351 4642 5439
rect 4700 5351 4900 5439
rect 4958 5401 5158 5439
rect 4958 5367 5007 5401
rect 5041 5367 5075 5401
rect 5109 5367 5158 5401
rect 4958 5351 5158 5367
rect 5216 5401 5416 5439
rect 5216 5367 5265 5401
rect 5299 5367 5333 5401
rect 5367 5367 5416 5401
rect 5216 5351 5416 5367
rect 5474 5351 5674 5439
rect 5732 5351 5932 5439
rect 5990 5401 6190 5439
rect 5990 5367 6039 5401
rect 6073 5367 6107 5401
rect 6141 5367 6190 5401
rect 5990 5351 6190 5367
rect 3668 5293 3868 5309
rect 3668 5259 3717 5293
rect 3751 5259 3785 5293
rect 3819 5259 3868 5293
rect 3668 5221 3868 5259
rect 3926 5293 4126 5309
rect 3926 5259 3975 5293
rect 4009 5259 4043 5293
rect 4077 5259 4126 5293
rect 3926 5221 4126 5259
rect 4184 5293 4384 5309
rect 4184 5259 4233 5293
rect 4267 5259 4301 5293
rect 4335 5259 4384 5293
rect 4184 5221 4384 5259
rect 4442 5221 4642 5309
rect 4700 5221 4900 5309
rect 4958 5293 5158 5309
rect 4958 5259 5007 5293
rect 5041 5259 5075 5293
rect 5109 5259 5158 5293
rect 4958 5221 5158 5259
rect 5216 5293 5416 5309
rect 5216 5259 5265 5293
rect 5299 5259 5333 5293
rect 5367 5259 5416 5293
rect 5216 5221 5416 5259
rect 5474 5221 5674 5309
rect 5732 5221 5932 5309
rect 5990 5293 6190 5309
rect 5990 5259 6039 5293
rect 6073 5259 6107 5293
rect 6141 5259 6190 5293
rect 5990 5221 6190 5259
rect 3668 4983 3868 5021
rect 3668 4949 3717 4983
rect 3751 4949 3785 4983
rect 3819 4949 3868 4983
rect 3668 4933 3868 4949
rect 3926 4933 4126 5021
rect 4184 4933 4384 5021
rect 4442 4983 4642 5021
rect 4442 4949 4491 4983
rect 4525 4949 4559 4983
rect 4593 4949 4642 4983
rect 4442 4933 4642 4949
rect 4700 4983 4900 5021
rect 4700 4949 4749 4983
rect 4783 4949 4817 4983
rect 4851 4949 4900 4983
rect 4700 4933 4900 4949
rect 4958 4933 5158 5021
rect 5216 4933 5416 5021
rect 5474 4983 5674 5021
rect 5474 4949 5523 4983
rect 5557 4949 5591 4983
rect 5625 4949 5674 4983
rect 5474 4933 5674 4949
rect 5732 4983 5932 5021
rect 5732 4949 5781 4983
rect 5815 4949 5849 4983
rect 5883 4949 5932 4983
rect 5732 4933 5932 4949
rect 5990 4983 6190 5021
rect 5990 4949 6039 4983
rect 6073 4949 6107 4983
rect 6141 4949 6190 4983
rect 5990 4933 6190 4949
rect 3668 4875 3868 4891
rect 3668 4841 3717 4875
rect 3751 4841 3785 4875
rect 3819 4841 3868 4875
rect 3668 4803 3868 4841
rect 3926 4803 4126 4891
rect 4184 4803 4384 4891
rect 4442 4875 4642 4891
rect 4442 4841 4491 4875
rect 4525 4841 4559 4875
rect 4593 4841 4642 4875
rect 4442 4803 4642 4841
rect 4700 4875 4900 4891
rect 4700 4841 4749 4875
rect 4783 4841 4817 4875
rect 4851 4841 4900 4875
rect 4700 4803 4900 4841
rect 4958 4803 5158 4891
rect 5216 4803 5416 4891
rect 5474 4875 5674 4891
rect 5474 4841 5523 4875
rect 5557 4841 5591 4875
rect 5625 4841 5674 4875
rect 5474 4803 5674 4841
rect 5732 4875 5932 4891
rect 5732 4841 5781 4875
rect 5815 4841 5849 4875
rect 5883 4841 5932 4875
rect 5732 4803 5932 4841
rect 5990 4875 6190 4891
rect 5990 4841 6039 4875
rect 6073 4841 6107 4875
rect 6141 4841 6190 4875
rect 5990 4803 6190 4841
rect 3668 4565 3868 4603
rect 3668 4531 3717 4565
rect 3751 4531 3785 4565
rect 3819 4531 3868 4565
rect 3668 4515 3868 4531
rect 3926 4565 4126 4603
rect 3926 4531 3975 4565
rect 4009 4531 4043 4565
rect 4077 4531 4126 4565
rect 3926 4515 4126 4531
rect 4184 4565 4384 4603
rect 4184 4531 4233 4565
rect 4267 4531 4301 4565
rect 4335 4531 4384 4565
rect 4184 4515 4384 4531
rect 4442 4515 4642 4603
rect 4700 4515 4900 4603
rect 4958 4565 5158 4603
rect 4958 4531 5007 4565
rect 5041 4531 5075 4565
rect 5109 4531 5158 4565
rect 4958 4515 5158 4531
rect 5216 4565 5416 4603
rect 5216 4531 5265 4565
rect 5299 4531 5333 4565
rect 5367 4531 5416 4565
rect 5216 4515 5416 4531
rect 5474 4515 5674 4603
rect 5732 4515 5932 4603
rect 5990 4565 6190 4603
rect 5990 4531 6039 4565
rect 6073 4531 6107 4565
rect 6141 4531 6190 4565
rect 5990 4515 6190 4531
rect 3668 4457 3868 4473
rect 3668 4423 3717 4457
rect 3751 4423 3785 4457
rect 3819 4423 3868 4457
rect 3668 4385 3868 4423
rect 3926 4457 4126 4473
rect 3926 4423 3975 4457
rect 4009 4423 4043 4457
rect 4077 4423 4126 4457
rect 3926 4385 4126 4423
rect 4184 4457 4384 4473
rect 4184 4423 4233 4457
rect 4267 4423 4301 4457
rect 4335 4423 4384 4457
rect 4184 4385 4384 4423
rect 4442 4457 4642 4473
rect 4442 4423 4491 4457
rect 4525 4423 4559 4457
rect 4593 4423 4642 4457
rect 4442 4385 4642 4423
rect 4700 4457 4900 4473
rect 4700 4423 4749 4457
rect 4783 4423 4817 4457
rect 4851 4423 4900 4457
rect 4700 4385 4900 4423
rect 4958 4457 5158 4473
rect 4958 4423 5007 4457
rect 5041 4423 5075 4457
rect 5109 4423 5158 4457
rect 4958 4385 5158 4423
rect 5216 4457 5416 4473
rect 5216 4423 5265 4457
rect 5299 4423 5333 4457
rect 5367 4423 5416 4457
rect 5216 4385 5416 4423
rect 5474 4457 5674 4473
rect 5474 4423 5523 4457
rect 5557 4423 5591 4457
rect 5625 4423 5674 4457
rect 5474 4385 5674 4423
rect 5732 4457 5932 4473
rect 5732 4423 5781 4457
rect 5815 4423 5849 4457
rect 5883 4423 5932 4457
rect 5732 4385 5932 4423
rect 5990 4457 6190 4473
rect 5990 4423 6039 4457
rect 6073 4423 6107 4457
rect 6141 4423 6190 4457
rect 5990 4385 6190 4423
rect 3668 4147 3868 4185
rect 3668 4113 3717 4147
rect 3751 4113 3785 4147
rect 3819 4113 3868 4147
rect 3668 4097 3868 4113
rect 3926 4097 4126 4185
rect 4184 4097 4384 4185
rect 4442 4097 4642 4185
rect 4700 4097 4900 4185
rect 4958 4097 5158 4185
rect 5216 4097 5416 4185
rect 5474 4097 5674 4185
rect 5732 4097 5932 4185
rect 5990 4147 6190 4185
rect 5990 4113 6039 4147
rect 6073 4113 6107 4147
rect 6141 4113 6190 4147
rect 5990 4097 6190 4113
rect 8404 6972 8604 6988
rect 8404 6938 8453 6972
rect 8487 6938 8521 6972
rect 8555 6938 8604 6972
rect 8404 6900 8604 6938
rect 8662 6972 8862 6988
rect 8662 6938 8711 6972
rect 8745 6938 8779 6972
rect 8813 6938 8862 6972
rect 8662 6900 8862 6938
rect 8920 6972 9120 6988
rect 8920 6938 8969 6972
rect 9003 6938 9037 6972
rect 9071 6938 9120 6972
rect 8920 6900 9120 6938
rect 9178 6972 9378 6988
rect 9178 6938 9227 6972
rect 9261 6938 9295 6972
rect 9329 6938 9378 6972
rect 9178 6900 9378 6938
rect 9436 6972 9636 6988
rect 9436 6938 9485 6972
rect 9519 6938 9553 6972
rect 9587 6938 9636 6972
rect 9436 6900 9636 6938
rect 9694 6972 9894 6988
rect 9694 6938 9743 6972
rect 9777 6938 9811 6972
rect 9845 6938 9894 6972
rect 9694 6900 9894 6938
rect 8404 6662 8604 6700
rect 8404 6628 8453 6662
rect 8487 6628 8521 6662
rect 8555 6628 8604 6662
rect 8404 6612 8604 6628
rect 8662 6612 8862 6700
rect 8920 6612 9120 6700
rect 9178 6612 9378 6700
rect 9436 6612 9636 6700
rect 9694 6662 9894 6700
rect 9694 6628 9743 6662
rect 9777 6628 9811 6662
rect 9845 6628 9894 6662
rect 9694 6612 9894 6628
rect 8404 6554 8604 6570
rect 8404 6520 8453 6554
rect 8487 6520 8521 6554
rect 8555 6520 8604 6554
rect 8404 6482 8604 6520
rect 8662 6554 8862 6570
rect 8662 6520 8711 6554
rect 8745 6520 8779 6554
rect 8813 6520 8862 6554
rect 8662 6482 8862 6520
rect 8920 6554 9120 6570
rect 8920 6520 8969 6554
rect 9003 6520 9037 6554
rect 9071 6520 9120 6554
rect 8920 6482 9120 6520
rect 9178 6554 9378 6570
rect 9178 6520 9227 6554
rect 9261 6520 9295 6554
rect 9329 6520 9378 6554
rect 9178 6482 9378 6520
rect 9436 6554 9636 6570
rect 9436 6520 9485 6554
rect 9519 6520 9553 6554
rect 9587 6520 9636 6554
rect 9436 6482 9636 6520
rect 9694 6554 9894 6570
rect 9694 6520 9743 6554
rect 9777 6520 9811 6554
rect 9845 6520 9894 6554
rect 9694 6482 9894 6520
rect 8404 6244 8604 6282
rect 8404 6210 8453 6244
rect 8487 6210 8521 6244
rect 8555 6210 8604 6244
rect 8404 6194 8604 6210
rect 8662 6194 8862 6282
rect 8920 6194 9120 6282
rect 9178 6194 9378 6282
rect 9436 6194 9636 6282
rect 9694 6244 9894 6282
rect 9694 6210 9743 6244
rect 9777 6210 9811 6244
rect 9845 6210 9894 6244
rect 9694 6194 9894 6210
rect 8404 6136 8604 6152
rect 8404 6102 8453 6136
rect 8487 6102 8521 6136
rect 8555 6102 8604 6136
rect 8404 6064 8604 6102
rect 8662 6136 8862 6152
rect 8662 6102 8711 6136
rect 8745 6102 8779 6136
rect 8813 6102 8862 6136
rect 8662 6064 8862 6102
rect 8920 6136 9120 6152
rect 8920 6102 8969 6136
rect 9003 6102 9037 6136
rect 9071 6102 9120 6136
rect 8920 6064 9120 6102
rect 9178 6136 9378 6152
rect 9178 6102 9227 6136
rect 9261 6102 9295 6136
rect 9329 6102 9378 6136
rect 9178 6064 9378 6102
rect 9436 6136 9636 6152
rect 9436 6102 9485 6136
rect 9519 6102 9553 6136
rect 9587 6102 9636 6136
rect 9436 6064 9636 6102
rect 9694 6136 9894 6152
rect 9694 6102 9743 6136
rect 9777 6102 9811 6136
rect 9845 6102 9894 6136
rect 9694 6064 9894 6102
rect 8404 5826 8604 5864
rect 8404 5792 8453 5826
rect 8487 5792 8521 5826
rect 8555 5792 8604 5826
rect 8404 5776 8604 5792
rect 8662 5776 8862 5864
rect 8920 5776 9120 5864
rect 9178 5776 9378 5864
rect 9436 5776 9636 5864
rect 9694 5826 9894 5864
rect 9694 5792 9743 5826
rect 9777 5792 9811 5826
rect 9845 5792 9894 5826
rect 9694 5776 9894 5792
rect 8404 5718 8604 5734
rect 8404 5684 8453 5718
rect 8487 5684 8521 5718
rect 8555 5684 8604 5718
rect 8404 5646 8604 5684
rect 8662 5718 8862 5734
rect 8662 5684 8711 5718
rect 8745 5684 8779 5718
rect 8813 5684 8862 5718
rect 8662 5646 8862 5684
rect 8920 5718 9120 5734
rect 8920 5684 8969 5718
rect 9003 5684 9037 5718
rect 9071 5684 9120 5718
rect 8920 5646 9120 5684
rect 9178 5718 9378 5734
rect 9178 5684 9227 5718
rect 9261 5684 9295 5718
rect 9329 5684 9378 5718
rect 9178 5646 9378 5684
rect 9436 5718 9636 5734
rect 9436 5684 9485 5718
rect 9519 5684 9553 5718
rect 9587 5684 9636 5718
rect 9436 5646 9636 5684
rect 9694 5718 9894 5734
rect 9694 5684 9743 5718
rect 9777 5684 9811 5718
rect 9845 5684 9894 5718
rect 9694 5646 9894 5684
rect 8404 5408 8604 5446
rect 8404 5374 8453 5408
rect 8487 5374 8521 5408
rect 8555 5374 8604 5408
rect 8404 5358 8604 5374
rect 8662 5358 8862 5446
rect 8920 5358 9120 5446
rect 9178 5358 9378 5446
rect 9436 5358 9636 5446
rect 9694 5408 9894 5446
rect 9694 5374 9743 5408
rect 9777 5374 9811 5408
rect 9845 5374 9894 5408
rect 9694 5358 9894 5374
rect 8404 5300 8604 5316
rect 8404 5266 8453 5300
rect 8487 5266 8521 5300
rect 8555 5266 8604 5300
rect 8404 5228 8604 5266
rect 8662 5300 8862 5316
rect 8662 5266 8711 5300
rect 8745 5266 8779 5300
rect 8813 5266 8862 5300
rect 8662 5228 8862 5266
rect 8920 5300 9120 5316
rect 8920 5266 8969 5300
rect 9003 5266 9037 5300
rect 9071 5266 9120 5300
rect 8920 5228 9120 5266
rect 9178 5300 9378 5316
rect 9178 5266 9227 5300
rect 9261 5266 9295 5300
rect 9329 5266 9378 5300
rect 9178 5228 9378 5266
rect 9436 5300 9636 5316
rect 9436 5266 9485 5300
rect 9519 5266 9553 5300
rect 9587 5266 9636 5300
rect 9436 5228 9636 5266
rect 9694 5300 9894 5316
rect 9694 5266 9743 5300
rect 9777 5266 9811 5300
rect 9845 5266 9894 5300
rect 9694 5228 9894 5266
rect 8404 4990 8604 5028
rect 8404 4956 8453 4990
rect 8487 4956 8521 4990
rect 8555 4956 8604 4990
rect 8404 4940 8604 4956
rect 8662 4940 8862 5028
rect 8920 4940 9120 5028
rect 9178 4940 9378 5028
rect 9436 4940 9636 5028
rect 9694 4990 9894 5028
rect 9694 4956 9743 4990
rect 9777 4956 9811 4990
rect 9845 4956 9894 4990
rect 9694 4940 9894 4956
rect 8404 4882 8604 4898
rect 8404 4848 8453 4882
rect 8487 4848 8521 4882
rect 8555 4848 8604 4882
rect 8404 4810 8604 4848
rect 8662 4882 8862 4898
rect 8662 4848 8711 4882
rect 8745 4848 8779 4882
rect 8813 4848 8862 4882
rect 8662 4810 8862 4848
rect 8920 4882 9120 4898
rect 8920 4848 8969 4882
rect 9003 4848 9037 4882
rect 9071 4848 9120 4882
rect 8920 4810 9120 4848
rect 9178 4882 9378 4898
rect 9178 4848 9227 4882
rect 9261 4848 9295 4882
rect 9329 4848 9378 4882
rect 9178 4810 9378 4848
rect 9436 4882 9636 4898
rect 9436 4848 9485 4882
rect 9519 4848 9553 4882
rect 9587 4848 9636 4882
rect 9436 4810 9636 4848
rect 9694 4882 9894 4898
rect 9694 4848 9743 4882
rect 9777 4848 9811 4882
rect 9845 4848 9894 4882
rect 9694 4810 9894 4848
rect 8404 4572 8604 4610
rect 8404 4538 8453 4572
rect 8487 4538 8521 4572
rect 8555 4538 8604 4572
rect 8404 4522 8604 4538
rect 8662 4522 8862 4610
rect 8920 4522 9120 4610
rect 9178 4522 9378 4610
rect 9436 4522 9636 4610
rect 9694 4572 9894 4610
rect 9694 4538 9743 4572
rect 9777 4538 9811 4572
rect 9845 4538 9894 4572
rect 9694 4522 9894 4538
rect 8404 4464 8604 4480
rect 8404 4430 8453 4464
rect 8487 4430 8521 4464
rect 8555 4430 8604 4464
rect 8404 4392 8604 4430
rect 8662 4464 8862 4480
rect 8662 4430 8711 4464
rect 8745 4430 8779 4464
rect 8813 4430 8862 4464
rect 8662 4392 8862 4430
rect 8920 4464 9120 4480
rect 8920 4430 8969 4464
rect 9003 4430 9037 4464
rect 9071 4430 9120 4464
rect 8920 4392 9120 4430
rect 9178 4464 9378 4480
rect 9178 4430 9227 4464
rect 9261 4430 9295 4464
rect 9329 4430 9378 4464
rect 9178 4392 9378 4430
rect 9436 4464 9636 4480
rect 9436 4430 9485 4464
rect 9519 4430 9553 4464
rect 9587 4430 9636 4464
rect 9436 4392 9636 4430
rect 9694 4464 9894 4480
rect 9694 4430 9743 4464
rect 9777 4430 9811 4464
rect 9845 4430 9894 4464
rect 9694 4392 9894 4430
rect 8404 4154 8604 4192
rect 8404 4120 8453 4154
rect 8487 4120 8521 4154
rect 8555 4120 8604 4154
rect 8404 4104 8604 4120
rect 8662 4104 8862 4192
rect 8920 4104 9120 4192
rect 9178 4104 9378 4192
rect 9436 4104 9636 4192
rect 9694 4154 9894 4192
rect 9694 4120 9743 4154
rect 9777 4120 9811 4154
rect 9845 4120 9894 4154
rect 9694 4104 9894 4120
rect -2162 3950 -1962 3988
rect -2162 3916 -2113 3950
rect -2079 3916 -2045 3950
rect -2011 3916 -1962 3950
rect -2162 3900 -1962 3916
rect -1904 3900 -1704 3988
rect -1646 3900 -1446 3988
rect -1388 3900 -1188 3988
rect -1130 3900 -930 3988
rect -872 3900 -672 3988
rect -614 3900 -414 3988
rect -356 3900 -156 3988
rect -98 3900 102 3988
rect 160 3900 360 3988
rect 418 3900 618 3988
rect 676 3900 876 3988
rect 934 3900 1134 3988
rect 1192 3950 1392 3988
rect 1192 3916 1241 3950
rect 1275 3916 1309 3950
rect 1343 3916 1392 3950
rect 1192 3900 1392 3916
<< polycont >>
rect 3178 10737 3212 10771
rect 3246 10737 3280 10771
rect 3436 10737 3470 10771
rect 3504 10737 3538 10771
rect 3694 10737 3728 10771
rect 3762 10737 3796 10771
rect 4468 10737 4502 10771
rect 4536 10737 4570 10771
rect 4726 10737 4760 10771
rect 4794 10737 4828 10771
rect 4984 10737 5018 10771
rect 5052 10737 5086 10771
rect -1144 10527 -1110 10561
rect -1076 10527 -1042 10561
rect 146 10527 180 10561
rect 214 10527 248 10561
rect -1144 10199 -1110 10233
rect -1076 10199 -1042 10233
rect -886 10199 -852 10233
rect -818 10199 -784 10233
rect -628 10199 -594 10233
rect -560 10199 -526 10233
rect -370 10199 -336 10233
rect -302 10199 -268 10233
rect -112 10199 -78 10233
rect -44 10199 -10 10233
rect 146 10199 180 10233
rect 214 10199 248 10233
rect -1144 10091 -1110 10125
rect -1076 10091 -1042 10125
rect -886 10091 -852 10125
rect -818 10091 -784 10125
rect -628 10091 -594 10125
rect -560 10091 -526 10125
rect -370 10091 -336 10125
rect -302 10091 -268 10125
rect -112 10091 -78 10125
rect -44 10091 -10 10125
rect 146 10091 180 10125
rect 214 10091 248 10125
rect -1144 9763 -1110 9797
rect -1076 9763 -1042 9797
rect 146 9763 180 9797
rect 214 9763 248 9797
rect -1144 9655 -1110 9689
rect -1076 9655 -1042 9689
rect 146 9655 180 9689
rect 214 9655 248 9689
rect -1144 9327 -1110 9361
rect -1076 9327 -1042 9361
rect -886 9327 -852 9361
rect -818 9327 -784 9361
rect -628 9327 -594 9361
rect -560 9327 -526 9361
rect -370 9327 -336 9361
rect -302 9327 -268 9361
rect -112 9327 -78 9361
rect -44 9327 -10 9361
rect 146 9327 180 9361
rect 214 9327 248 9361
rect -1144 9219 -1110 9253
rect -1076 9219 -1042 9253
rect -886 9219 -852 9253
rect -818 9219 -784 9253
rect -628 9219 -594 9253
rect -560 9219 -526 9253
rect -370 9219 -336 9253
rect -302 9219 -268 9253
rect -112 9219 -78 9253
rect -44 9219 -10 9253
rect 146 9219 180 9253
rect 214 9219 248 9253
rect -1144 8891 -1110 8925
rect -1076 8891 -1042 8925
rect 146 8891 180 8925
rect 214 8891 248 8925
rect 3178 10427 3212 10461
rect 3246 10427 3280 10461
rect 3952 10427 3986 10461
rect 4020 10427 4054 10461
rect 4210 10427 4244 10461
rect 4278 10427 4312 10461
rect 4984 10424 5018 10458
rect 5052 10424 5086 10458
rect 3178 10319 3212 10353
rect 3246 10319 3280 10353
rect 3952 10319 3986 10353
rect 4020 10319 4054 10353
rect 4210 10319 4244 10353
rect 4278 10319 4312 10353
rect 4984 10319 5018 10353
rect 5052 10319 5086 10353
rect 3178 10009 3212 10043
rect 3246 10009 3280 10043
rect 3436 10009 3470 10043
rect 3504 10009 3538 10043
rect 3694 10009 3728 10043
rect 3762 10009 3796 10043
rect 4468 10009 4502 10043
rect 4536 10009 4570 10043
rect 4726 10009 4760 10043
rect 4794 10009 4828 10043
rect 4984 10009 5018 10043
rect 5052 10009 5086 10043
rect 3178 9901 3212 9935
rect 3246 9901 3280 9935
rect 3436 9901 3470 9935
rect 3504 9901 3538 9935
rect 3694 9901 3728 9935
rect 3762 9901 3796 9935
rect 4468 9901 4502 9935
rect 4536 9901 4570 9935
rect 4726 9901 4760 9935
rect 4794 9901 4828 9935
rect 4984 9901 5018 9935
rect 5052 9901 5086 9935
rect 3178 9591 3212 9625
rect 3246 9591 3280 9625
rect 3952 9591 3986 9625
rect 4020 9591 4054 9625
rect 4210 9591 4244 9625
rect 4278 9591 4312 9625
rect 4984 9588 5018 9622
rect 5052 9588 5086 9622
rect 3178 9483 3212 9517
rect 3246 9483 3280 9517
rect 3952 9483 3986 9517
rect 4020 9483 4054 9517
rect 4210 9483 4244 9517
rect 4278 9483 4312 9517
rect 4984 9483 5018 9517
rect 5052 9483 5086 9517
rect 3178 9173 3212 9207
rect 3246 9173 3280 9207
rect 3436 9173 3470 9207
rect 3504 9173 3538 9207
rect 3694 9173 3728 9207
rect 3762 9173 3796 9207
rect 4468 9173 4502 9207
rect 4536 9173 4570 9207
rect 4726 9173 4760 9207
rect 4794 9173 4828 9207
rect 4984 9170 5018 9204
rect 5052 9170 5086 9204
rect 3178 9061 3212 9095
rect 3246 9061 3280 9095
rect 3436 9061 3470 9095
rect 3504 9061 3538 9095
rect 3694 9061 3728 9095
rect 3762 9061 3796 9095
rect 4468 9061 4502 9095
rect 4536 9061 4570 9095
rect 4726 9061 4760 9095
rect 4794 9061 4828 9095
rect 4984 9061 5018 9095
rect 5052 9061 5086 9095
rect 3178 8751 3212 8785
rect 3246 8751 3280 8785
rect 3952 8751 3986 8785
rect 4020 8751 4054 8785
rect 4210 8751 4244 8785
rect 4278 8751 4312 8785
rect 4984 8748 5018 8782
rect 5052 8748 5086 8782
rect 3178 8639 3212 8673
rect 3246 8639 3280 8673
rect 3952 8639 3986 8673
rect 4020 8639 4054 8673
rect 4210 8639 4244 8673
rect 4278 8639 4312 8673
rect 4984 8639 5018 8673
rect 5052 8639 5086 8673
rect 3178 8329 3212 8363
rect 3246 8329 3280 8363
rect 3436 8329 3470 8363
rect 3504 8329 3538 8363
rect 3694 8329 3728 8363
rect 3762 8329 3796 8363
rect 4468 8329 4502 8363
rect 4536 8329 4570 8363
rect 4726 8329 4760 8363
rect 4794 8329 4828 8363
rect 4984 8329 5018 8363
rect 5052 8329 5086 8363
rect 7104 10845 7138 10879
rect 7172 10845 7206 10879
rect 8394 10845 8428 10879
rect 8462 10845 8496 10879
rect 7104 10517 7138 10551
rect 7172 10517 7206 10551
rect 7362 10517 7396 10551
rect 7430 10517 7464 10551
rect 7620 10517 7654 10551
rect 7688 10517 7722 10551
rect 7878 10517 7912 10551
rect 7946 10517 7980 10551
rect 8136 10517 8170 10551
rect 8204 10517 8238 10551
rect 8394 10517 8428 10551
rect 8462 10517 8496 10551
rect 7104 10409 7138 10443
rect 7172 10409 7206 10443
rect 7362 10409 7396 10443
rect 7430 10409 7464 10443
rect 7620 10409 7654 10443
rect 7688 10409 7722 10443
rect 7878 10409 7912 10443
rect 7946 10409 7980 10443
rect 8136 10409 8170 10443
rect 8204 10409 8238 10443
rect 8394 10409 8428 10443
rect 8462 10409 8496 10443
rect 7104 10081 7138 10115
rect 7172 10081 7206 10115
rect 8394 10081 8428 10115
rect 8462 10081 8496 10115
rect 7104 9973 7138 10007
rect 7172 9973 7206 10007
rect 8394 9973 8428 10007
rect 8462 9973 8496 10007
rect 7104 9645 7138 9679
rect 7172 9645 7206 9679
rect 7362 9645 7396 9679
rect 7430 9645 7464 9679
rect 7620 9645 7654 9679
rect 7688 9645 7722 9679
rect 7878 9645 7912 9679
rect 7946 9645 7980 9679
rect 8136 9645 8170 9679
rect 8204 9645 8238 9679
rect 8394 9645 8428 9679
rect 8462 9645 8496 9679
rect 7104 9537 7138 9571
rect 7172 9537 7206 9571
rect 7362 9537 7396 9571
rect 7430 9537 7464 9571
rect 7620 9537 7654 9571
rect 7688 9537 7722 9571
rect 7878 9537 7912 9571
rect 7946 9537 7980 9571
rect 8136 9537 8170 9571
rect 8204 9537 8238 9571
rect 8394 9537 8428 9571
rect 8462 9537 8496 9571
rect 7104 9209 7138 9243
rect 7172 9209 7206 9243
rect 8394 9209 8428 9243
rect 8462 9209 8496 9243
rect 7104 9101 7138 9135
rect 7172 9101 7206 9135
rect 8394 9101 8428 9135
rect 8462 9101 8496 9135
rect 7104 8773 7138 8807
rect 7172 8773 7206 8807
rect 7362 8773 7396 8807
rect 7430 8773 7464 8807
rect 7620 8773 7654 8807
rect 7688 8773 7722 8807
rect 7878 8773 7912 8807
rect 7946 8773 7980 8807
rect 8136 8773 8170 8807
rect 8204 8773 8238 8807
rect 8394 8773 8428 8807
rect 8462 8773 8496 8807
rect 7104 8665 7138 8699
rect 7172 8665 7206 8699
rect 7362 8665 7396 8699
rect 7430 8665 7464 8699
rect 7620 8665 7654 8699
rect 7688 8665 7722 8699
rect 7878 8665 7912 8699
rect 7946 8665 7980 8699
rect 8136 8665 8170 8699
rect 8204 8665 8238 8699
rect 8394 8665 8428 8699
rect 8462 8665 8496 8699
rect 7104 8337 7138 8371
rect 7172 8337 7206 8371
rect 8394 8337 8428 8371
rect 8462 8337 8496 8371
rect 7104 8229 7138 8263
rect 7172 8229 7206 8263
rect 7362 8229 7396 8263
rect 7430 8229 7464 8263
rect 7620 8229 7654 8263
rect 7688 8229 7722 8263
rect 7878 8229 7912 8263
rect 7946 8229 7980 8263
rect 8136 8229 8170 8263
rect 8204 8229 8238 8263
rect 8394 8229 8428 8263
rect 8462 8229 8496 8263
rect -2113 7988 -2079 8022
rect -2045 7988 -2011 8022
rect -1855 7988 -1821 8022
rect -1787 7988 -1753 8022
rect -1597 7988 -1563 8022
rect -1529 7988 -1495 8022
rect -1339 7988 -1305 8022
rect -1271 7988 -1237 8022
rect -1081 7988 -1047 8022
rect -1013 7988 -979 8022
rect -823 7988 -789 8022
rect -755 7988 -721 8022
rect -565 7988 -531 8022
rect -497 7988 -463 8022
rect -307 7988 -273 8022
rect -239 7988 -205 8022
rect -49 7988 -15 8022
rect 19 7988 53 8022
rect 209 7988 243 8022
rect 277 7988 311 8022
rect 467 7988 501 8022
rect 535 7988 569 8022
rect 725 7988 759 8022
rect 793 7988 827 8022
rect 983 7988 1017 8022
rect 1051 7988 1085 8022
rect 1241 7988 1275 8022
rect 1309 7988 1343 8022
rect 7104 7901 7138 7935
rect 7172 7901 7206 7935
rect 8394 7901 8428 7935
rect 8462 7901 8496 7935
rect -2113 7678 -2079 7712
rect -2045 7678 -2011 7712
rect 1241 7678 1275 7712
rect 1309 7678 1343 7712
rect -2113 7570 -2079 7604
rect -2045 7570 -2011 7604
rect -1855 7570 -1821 7604
rect -1787 7570 -1753 7604
rect -1597 7570 -1563 7604
rect -1529 7570 -1495 7604
rect -1339 7570 -1305 7604
rect -1271 7570 -1237 7604
rect -1081 7570 -1047 7604
rect -1013 7570 -979 7604
rect -307 7570 -273 7604
rect -239 7570 -205 7604
rect -49 7570 -15 7604
rect 19 7570 53 7604
rect 725 7570 759 7604
rect 793 7570 827 7604
rect 983 7570 1017 7604
rect 1051 7570 1085 7604
rect 1241 7570 1275 7604
rect 1309 7570 1343 7604
rect -2113 7260 -2079 7294
rect -2045 7260 -2011 7294
rect -823 7260 -789 7294
rect -755 7260 -721 7294
rect -565 7260 -531 7294
rect -497 7260 -463 7294
rect 209 7260 243 7294
rect 277 7260 311 7294
rect 467 7260 501 7294
rect 535 7260 569 7294
rect 1241 7260 1275 7294
rect 1309 7260 1343 7294
rect -2113 7152 -2079 7186
rect -2045 7152 -2011 7186
rect -1855 7152 -1821 7186
rect -1787 7152 -1753 7186
rect -1597 7152 -1563 7186
rect -1529 7152 -1495 7186
rect -823 7152 -789 7186
rect -755 7152 -721 7186
rect -565 7152 -531 7186
rect -497 7152 -463 7186
rect 209 7152 243 7186
rect 277 7152 311 7186
rect 467 7152 501 7186
rect 535 7152 569 7186
rect 1241 7152 1275 7186
rect 1309 7152 1343 7186
rect -2113 6842 -2079 6876
rect -2045 6842 -2011 6876
rect -1339 6842 -1305 6876
rect -1271 6842 -1237 6876
rect -1081 6842 -1047 6876
rect -1013 6842 -979 6876
rect -307 6842 -273 6876
rect -239 6842 -205 6876
rect -49 6842 -15 6876
rect 19 6842 53 6876
rect 725 6842 759 6876
rect 793 6842 827 6876
rect 983 6842 1017 6876
rect 1051 6842 1085 6876
rect 1241 6842 1275 6876
rect 1309 6842 1343 6876
rect -2113 6734 -2079 6768
rect -2045 6734 -2011 6768
rect -1339 6734 -1305 6768
rect -1271 6734 -1237 6768
rect -1081 6734 -1047 6768
rect -1013 6734 -979 6768
rect -307 6734 -273 6768
rect -239 6734 -205 6768
rect -49 6734 -15 6768
rect 19 6734 53 6768
rect 725 6734 759 6768
rect 793 6734 827 6768
rect 983 6734 1017 6768
rect 1051 6734 1085 6768
rect 1241 6734 1275 6768
rect 1309 6734 1343 6768
rect -2113 6424 -2079 6458
rect -2045 6424 -2011 6458
rect -1855 6424 -1821 6458
rect -1787 6424 -1753 6458
rect -1597 6424 -1563 6458
rect -1529 6424 -1495 6458
rect -823 6424 -789 6458
rect -755 6424 -721 6458
rect -565 6424 -531 6458
rect -497 6424 -463 6458
rect 209 6424 243 6458
rect 277 6424 311 6458
rect 467 6424 501 6458
rect 535 6424 569 6458
rect 1241 6424 1275 6458
rect 1309 6424 1343 6458
rect -2113 6316 -2079 6350
rect -2045 6316 -2011 6350
rect -1855 6316 -1821 6350
rect -1787 6316 -1753 6350
rect -1597 6316 -1563 6350
rect -1529 6316 -1495 6350
rect -823 6316 -789 6350
rect -755 6316 -721 6350
rect -565 6316 -531 6350
rect -497 6316 -463 6350
rect 209 6316 243 6350
rect 277 6316 311 6350
rect 467 6316 501 6350
rect 535 6316 569 6350
rect 1241 6316 1275 6350
rect 1309 6316 1343 6350
rect -2113 6006 -2079 6040
rect -2045 6006 -2011 6040
rect -1339 6006 -1305 6040
rect -1271 6006 -1237 6040
rect -1081 6006 -1047 6040
rect -1013 6006 -979 6040
rect -307 6006 -273 6040
rect -239 6006 -205 6040
rect -49 6006 -15 6040
rect 19 6006 53 6040
rect 725 6006 759 6040
rect 793 6006 827 6040
rect 983 6006 1017 6040
rect 1051 6006 1085 6040
rect 1241 6006 1275 6040
rect 1309 6006 1343 6040
rect -2113 5898 -2079 5932
rect -2045 5898 -2011 5932
rect -1339 5898 -1305 5932
rect -1271 5898 -1237 5932
rect -1081 5898 -1047 5932
rect -1013 5898 -979 5932
rect -307 5898 -273 5932
rect -239 5898 -205 5932
rect -49 5898 -15 5932
rect 19 5898 53 5932
rect 725 5898 759 5932
rect 793 5898 827 5932
rect 983 5898 1017 5932
rect 1051 5898 1085 5932
rect 1241 5898 1275 5932
rect 1309 5898 1343 5932
rect -2113 5588 -2079 5622
rect -2045 5588 -2011 5622
rect -1855 5588 -1821 5622
rect -1787 5588 -1753 5622
rect -1597 5588 -1563 5622
rect -1529 5588 -1495 5622
rect -823 5588 -789 5622
rect -755 5588 -721 5622
rect -565 5588 -531 5622
rect -497 5588 -463 5622
rect 209 5588 243 5622
rect 277 5588 311 5622
rect 467 5588 501 5622
rect 535 5588 569 5622
rect 1241 5588 1275 5622
rect 1309 5588 1343 5622
rect -2113 5480 -2079 5514
rect -2045 5480 -2011 5514
rect -1855 5480 -1821 5514
rect -1787 5480 -1753 5514
rect -1597 5480 -1563 5514
rect -1529 5480 -1495 5514
rect -823 5480 -789 5514
rect -755 5480 -721 5514
rect -565 5480 -531 5514
rect -497 5480 -463 5514
rect 209 5480 243 5514
rect 277 5480 311 5514
rect 467 5480 501 5514
rect 535 5480 569 5514
rect 1241 5480 1275 5514
rect 1309 5480 1343 5514
rect -2113 5170 -2079 5204
rect -2045 5170 -2011 5204
rect -1339 5170 -1305 5204
rect -1271 5170 -1237 5204
rect -1081 5170 -1047 5204
rect -1013 5170 -979 5204
rect -307 5170 -273 5204
rect -239 5170 -205 5204
rect -49 5170 -15 5204
rect 19 5170 53 5204
rect 725 5170 759 5204
rect 793 5170 827 5204
rect 983 5170 1017 5204
rect 1051 5170 1085 5204
rect 1241 5170 1275 5204
rect 1309 5170 1343 5204
rect -2113 5062 -2079 5096
rect -2045 5062 -2011 5096
rect -1339 5062 -1305 5096
rect -1271 5062 -1237 5096
rect -1081 5062 -1047 5096
rect -1013 5062 -979 5096
rect -307 5062 -273 5096
rect -239 5062 -205 5096
rect -49 5062 -15 5096
rect 19 5062 53 5096
rect 725 5062 759 5096
rect 793 5062 827 5096
rect 983 5062 1017 5096
rect 1051 5062 1085 5096
rect 1241 5062 1275 5096
rect 1309 5062 1343 5096
rect -2113 4752 -2079 4786
rect -2045 4752 -2011 4786
rect -1855 4752 -1821 4786
rect -1787 4752 -1753 4786
rect -1597 4752 -1563 4786
rect -1529 4752 -1495 4786
rect -823 4752 -789 4786
rect -755 4752 -721 4786
rect -565 4752 -531 4786
rect -497 4752 -463 4786
rect 209 4752 243 4786
rect 277 4752 311 4786
rect 467 4752 501 4786
rect 535 4752 569 4786
rect 1241 4752 1275 4786
rect 1309 4752 1343 4786
rect -2113 4644 -2079 4678
rect -2045 4644 -2011 4678
rect -1855 4644 -1821 4678
rect -1787 4644 -1753 4678
rect -1597 4644 -1563 4678
rect -1529 4644 -1495 4678
rect -823 4644 -789 4678
rect -755 4644 -721 4678
rect -565 4644 -531 4678
rect -497 4644 -463 4678
rect 209 4644 243 4678
rect 277 4644 311 4678
rect 467 4644 501 4678
rect 535 4644 569 4678
rect 725 4644 759 4678
rect 793 4644 827 4678
rect 983 4644 1017 4678
rect 1051 4644 1085 4678
rect 1241 4644 1275 4678
rect 1309 4644 1343 4678
rect -2113 4334 -2079 4368
rect -2045 4334 -2011 4368
rect -1339 4334 -1305 4368
rect -1271 4334 -1237 4368
rect -1081 4334 -1047 4368
rect -1013 4334 -979 4368
rect -307 4334 -273 4368
rect -239 4334 -205 4368
rect -49 4334 -15 4368
rect 19 4334 53 4368
rect 1241 4334 1275 4368
rect 1309 4334 1343 4368
rect -2113 4226 -2079 4260
rect -2045 4226 -2011 4260
rect -1855 4226 -1821 4260
rect -1787 4226 -1753 4260
rect -1597 4226 -1563 4260
rect -1529 4226 -1495 4260
rect -1339 4226 -1305 4260
rect -1271 4226 -1237 4260
rect -1081 4226 -1047 4260
rect -1013 4226 -979 4260
rect -823 4226 -789 4260
rect -755 4226 -721 4260
rect -565 4226 -531 4260
rect -497 4226 -463 4260
rect -307 4226 -273 4260
rect -239 4226 -205 4260
rect -49 4226 -15 4260
rect 19 4226 53 4260
rect 209 4226 243 4260
rect 277 4226 311 4260
rect 467 4226 501 4260
rect 535 4226 569 4260
rect 725 4226 759 4260
rect 793 4226 827 4260
rect 983 4226 1017 4260
rect 1051 4226 1085 4260
rect 1241 4226 1275 4260
rect 1309 4226 1343 4260
rect 3717 7349 3751 7383
rect 3785 7349 3819 7383
rect 3975 7349 4009 7383
rect 4043 7349 4077 7383
rect 4233 7349 4267 7383
rect 4301 7349 4335 7383
rect 4491 7349 4525 7383
rect 4559 7349 4593 7383
rect 4749 7349 4783 7383
rect 4817 7349 4851 7383
rect 5007 7349 5041 7383
rect 5075 7349 5109 7383
rect 5265 7349 5299 7383
rect 5333 7349 5367 7383
rect 5523 7349 5557 7383
rect 5591 7349 5625 7383
rect 5781 7349 5815 7383
rect 5849 7349 5883 7383
rect 6039 7349 6073 7383
rect 6107 7349 6141 7383
rect 3717 7039 3751 7073
rect 3785 7039 3819 7073
rect 6039 7039 6073 7073
rect 6107 7039 6141 7073
rect 3717 6931 3751 6965
rect 3785 6931 3819 6965
rect 3975 6931 4009 6965
rect 4043 6931 4077 6965
rect 4233 6931 4267 6965
rect 4301 6931 4335 6965
rect 5007 6931 5041 6965
rect 5075 6931 5109 6965
rect 5265 6931 5299 6965
rect 5333 6931 5367 6965
rect 6039 6931 6073 6965
rect 6107 6931 6141 6965
rect 3717 6621 3751 6655
rect 3785 6621 3819 6655
rect 4491 6621 4525 6655
rect 4559 6621 4593 6655
rect 4749 6621 4783 6655
rect 4817 6621 4851 6655
rect 5523 6621 5557 6655
rect 5591 6621 5625 6655
rect 5781 6621 5815 6655
rect 5849 6621 5883 6655
rect 6039 6621 6073 6655
rect 6107 6621 6141 6655
rect 3717 6513 3751 6547
rect 3785 6513 3819 6547
rect 4491 6513 4525 6547
rect 4559 6513 4593 6547
rect 4749 6513 4783 6547
rect 4817 6513 4851 6547
rect 5523 6513 5557 6547
rect 5591 6513 5625 6547
rect 5781 6513 5815 6547
rect 5849 6513 5883 6547
rect 6039 6513 6073 6547
rect 6107 6513 6141 6547
rect 3717 6203 3751 6237
rect 3785 6203 3819 6237
rect 3975 6203 4009 6237
rect 4043 6203 4077 6237
rect 4233 6203 4267 6237
rect 4301 6203 4335 6237
rect 5007 6203 5041 6237
rect 5075 6203 5109 6237
rect 5265 6203 5299 6237
rect 5333 6203 5367 6237
rect 6039 6203 6073 6237
rect 6107 6203 6141 6237
rect 3717 6095 3751 6129
rect 3785 6095 3819 6129
rect 3975 6095 4009 6129
rect 4043 6095 4077 6129
rect 4233 6095 4267 6129
rect 4301 6095 4335 6129
rect 5007 6095 5041 6129
rect 5075 6095 5109 6129
rect 5265 6095 5299 6129
rect 5333 6095 5367 6129
rect 6039 6095 6073 6129
rect 6107 6095 6141 6129
rect 3717 5785 3751 5819
rect 3785 5785 3819 5819
rect 4491 5785 4525 5819
rect 4559 5785 4593 5819
rect 4749 5785 4783 5819
rect 4817 5785 4851 5819
rect 5523 5785 5557 5819
rect 5591 5785 5625 5819
rect 5781 5785 5815 5819
rect 5849 5785 5883 5819
rect 6039 5785 6073 5819
rect 6107 5785 6141 5819
rect 3717 5677 3751 5711
rect 3785 5677 3819 5711
rect 4491 5677 4525 5711
rect 4559 5677 4593 5711
rect 4749 5677 4783 5711
rect 4817 5677 4851 5711
rect 5523 5677 5557 5711
rect 5591 5677 5625 5711
rect 5781 5677 5815 5711
rect 5849 5677 5883 5711
rect 6039 5677 6073 5711
rect 6107 5677 6141 5711
rect 3717 5367 3751 5401
rect 3785 5367 3819 5401
rect 3975 5367 4009 5401
rect 4043 5367 4077 5401
rect 4233 5367 4267 5401
rect 4301 5367 4335 5401
rect 5007 5367 5041 5401
rect 5075 5367 5109 5401
rect 5265 5367 5299 5401
rect 5333 5367 5367 5401
rect 6039 5367 6073 5401
rect 6107 5367 6141 5401
rect 3717 5259 3751 5293
rect 3785 5259 3819 5293
rect 3975 5259 4009 5293
rect 4043 5259 4077 5293
rect 4233 5259 4267 5293
rect 4301 5259 4335 5293
rect 5007 5259 5041 5293
rect 5075 5259 5109 5293
rect 5265 5259 5299 5293
rect 5333 5259 5367 5293
rect 6039 5259 6073 5293
rect 6107 5259 6141 5293
rect 3717 4949 3751 4983
rect 3785 4949 3819 4983
rect 4491 4949 4525 4983
rect 4559 4949 4593 4983
rect 4749 4949 4783 4983
rect 4817 4949 4851 4983
rect 5523 4949 5557 4983
rect 5591 4949 5625 4983
rect 5781 4949 5815 4983
rect 5849 4949 5883 4983
rect 6039 4949 6073 4983
rect 6107 4949 6141 4983
rect 3717 4841 3751 4875
rect 3785 4841 3819 4875
rect 4491 4841 4525 4875
rect 4559 4841 4593 4875
rect 4749 4841 4783 4875
rect 4817 4841 4851 4875
rect 5523 4841 5557 4875
rect 5591 4841 5625 4875
rect 5781 4841 5815 4875
rect 5849 4841 5883 4875
rect 6039 4841 6073 4875
rect 6107 4841 6141 4875
rect 3717 4531 3751 4565
rect 3785 4531 3819 4565
rect 3975 4531 4009 4565
rect 4043 4531 4077 4565
rect 4233 4531 4267 4565
rect 4301 4531 4335 4565
rect 5007 4531 5041 4565
rect 5075 4531 5109 4565
rect 5265 4531 5299 4565
rect 5333 4531 5367 4565
rect 6039 4531 6073 4565
rect 6107 4531 6141 4565
rect 3717 4423 3751 4457
rect 3785 4423 3819 4457
rect 3975 4423 4009 4457
rect 4043 4423 4077 4457
rect 4233 4423 4267 4457
rect 4301 4423 4335 4457
rect 4491 4423 4525 4457
rect 4559 4423 4593 4457
rect 4749 4423 4783 4457
rect 4817 4423 4851 4457
rect 5007 4423 5041 4457
rect 5075 4423 5109 4457
rect 5265 4423 5299 4457
rect 5333 4423 5367 4457
rect 5523 4423 5557 4457
rect 5591 4423 5625 4457
rect 5781 4423 5815 4457
rect 5849 4423 5883 4457
rect 6039 4423 6073 4457
rect 6107 4423 6141 4457
rect 3717 4113 3751 4147
rect 3785 4113 3819 4147
rect 6039 4113 6073 4147
rect 6107 4113 6141 4147
rect 8453 6938 8487 6972
rect 8521 6938 8555 6972
rect 8711 6938 8745 6972
rect 8779 6938 8813 6972
rect 8969 6938 9003 6972
rect 9037 6938 9071 6972
rect 9227 6938 9261 6972
rect 9295 6938 9329 6972
rect 9485 6938 9519 6972
rect 9553 6938 9587 6972
rect 9743 6938 9777 6972
rect 9811 6938 9845 6972
rect 8453 6628 8487 6662
rect 8521 6628 8555 6662
rect 9743 6628 9777 6662
rect 9811 6628 9845 6662
rect 8453 6520 8487 6554
rect 8521 6520 8555 6554
rect 8711 6520 8745 6554
rect 8779 6520 8813 6554
rect 8969 6520 9003 6554
rect 9037 6520 9071 6554
rect 9227 6520 9261 6554
rect 9295 6520 9329 6554
rect 9485 6520 9519 6554
rect 9553 6520 9587 6554
rect 9743 6520 9777 6554
rect 9811 6520 9845 6554
rect 8453 6210 8487 6244
rect 8521 6210 8555 6244
rect 9743 6210 9777 6244
rect 9811 6210 9845 6244
rect 8453 6102 8487 6136
rect 8521 6102 8555 6136
rect 8711 6102 8745 6136
rect 8779 6102 8813 6136
rect 8969 6102 9003 6136
rect 9037 6102 9071 6136
rect 9227 6102 9261 6136
rect 9295 6102 9329 6136
rect 9485 6102 9519 6136
rect 9553 6102 9587 6136
rect 9743 6102 9777 6136
rect 9811 6102 9845 6136
rect 8453 5792 8487 5826
rect 8521 5792 8555 5826
rect 9743 5792 9777 5826
rect 9811 5792 9845 5826
rect 8453 5684 8487 5718
rect 8521 5684 8555 5718
rect 8711 5684 8745 5718
rect 8779 5684 8813 5718
rect 8969 5684 9003 5718
rect 9037 5684 9071 5718
rect 9227 5684 9261 5718
rect 9295 5684 9329 5718
rect 9485 5684 9519 5718
rect 9553 5684 9587 5718
rect 9743 5684 9777 5718
rect 9811 5684 9845 5718
rect 8453 5374 8487 5408
rect 8521 5374 8555 5408
rect 9743 5374 9777 5408
rect 9811 5374 9845 5408
rect 8453 5266 8487 5300
rect 8521 5266 8555 5300
rect 8711 5266 8745 5300
rect 8779 5266 8813 5300
rect 8969 5266 9003 5300
rect 9037 5266 9071 5300
rect 9227 5266 9261 5300
rect 9295 5266 9329 5300
rect 9485 5266 9519 5300
rect 9553 5266 9587 5300
rect 9743 5266 9777 5300
rect 9811 5266 9845 5300
rect 8453 4956 8487 4990
rect 8521 4956 8555 4990
rect 9743 4956 9777 4990
rect 9811 4956 9845 4990
rect 8453 4848 8487 4882
rect 8521 4848 8555 4882
rect 8711 4848 8745 4882
rect 8779 4848 8813 4882
rect 8969 4848 9003 4882
rect 9037 4848 9071 4882
rect 9227 4848 9261 4882
rect 9295 4848 9329 4882
rect 9485 4848 9519 4882
rect 9553 4848 9587 4882
rect 9743 4848 9777 4882
rect 9811 4848 9845 4882
rect 8453 4538 8487 4572
rect 8521 4538 8555 4572
rect 9743 4538 9777 4572
rect 9811 4538 9845 4572
rect 8453 4430 8487 4464
rect 8521 4430 8555 4464
rect 8711 4430 8745 4464
rect 8779 4430 8813 4464
rect 8969 4430 9003 4464
rect 9037 4430 9071 4464
rect 9227 4430 9261 4464
rect 9295 4430 9329 4464
rect 9485 4430 9519 4464
rect 9553 4430 9587 4464
rect 9743 4430 9777 4464
rect 9811 4430 9845 4464
rect 8453 4120 8487 4154
rect 8521 4120 8555 4154
rect 9743 4120 9777 4154
rect 9811 4120 9845 4154
rect -2113 3916 -2079 3950
rect -2045 3916 -2011 3950
rect 1241 3916 1275 3950
rect 1309 3916 1343 3950
<< locali >>
rect 6895 10947 7015 10981
rect 7049 10947 7083 10981
rect 7117 10947 7151 10981
rect 7185 10947 7219 10981
rect 7253 10947 7287 10981
rect 7321 10947 7355 10981
rect 7389 10947 7423 10981
rect 7457 10947 7491 10981
rect 7525 10947 7559 10981
rect 7593 10947 7627 10981
rect 7661 10947 7695 10981
rect 7729 10947 7763 10981
rect 7797 10947 7831 10981
rect 7865 10947 7899 10981
rect 7933 10947 7967 10981
rect 8001 10947 8035 10981
rect 8069 10947 8103 10981
rect 8137 10947 8171 10981
rect 8205 10947 8239 10981
rect 8273 10947 8299 10981
rect 8341 10947 8375 10981
rect 8409 10947 8443 10981
rect 8477 10947 8511 10981
rect 8545 10947 8579 10981
rect 8613 10947 8705 10981
rect 2969 10839 3089 10873
rect 3123 10839 3157 10873
rect 3191 10839 3225 10873
rect 3259 10839 3293 10873
rect 3327 10839 3361 10873
rect 3395 10839 3429 10873
rect 3463 10839 3497 10873
rect 3531 10839 3565 10873
rect 3599 10839 3633 10873
rect 3667 10839 3701 10873
rect 3735 10839 3769 10873
rect 3803 10839 3837 10873
rect 3871 10839 3905 10873
rect 3939 10839 3973 10873
rect 4007 10839 4041 10873
rect 4075 10839 4109 10873
rect 4143 10839 4177 10873
rect 4211 10839 4245 10873
rect 4279 10839 4313 10873
rect 4347 10839 4381 10873
rect 4415 10839 4449 10873
rect 4483 10839 4517 10873
rect 4551 10839 4585 10873
rect 4619 10839 4653 10873
rect 4687 10839 4721 10873
rect 4755 10839 4789 10873
rect 4823 10839 4857 10873
rect 4891 10839 4925 10873
rect 4959 10839 4993 10873
rect 5027 10839 5061 10873
rect 5095 10839 5129 10873
rect 5163 10839 5296 10873
rect 2969 10771 3003 10839
rect 5262 10771 5296 10839
rect 3129 10737 3176 10771
rect 3212 10737 3246 10771
rect 3282 10737 3329 10771
rect 3387 10737 3434 10771
rect 3470 10737 3504 10771
rect 3540 10737 3587 10771
rect 3645 10737 3692 10771
rect 3728 10737 3762 10771
rect 3798 10737 3845 10771
rect 4419 10737 4466 10771
rect 4502 10737 4536 10771
rect 4572 10737 4619 10771
rect 4677 10737 4724 10771
rect 4760 10737 4794 10771
rect 4830 10737 4877 10771
rect 4935 10737 4982 10771
rect 5018 10737 5052 10771
rect 5088 10737 5135 10771
rect 2969 10703 3003 10737
rect 5262 10703 5296 10737
rect -1353 10629 -1239 10663
rect -1199 10629 -1165 10663
rect -1131 10629 -1097 10663
rect -1063 10629 -1029 10663
rect -995 10629 -961 10663
rect -927 10629 -893 10663
rect -859 10629 -825 10663
rect -791 10629 -757 10663
rect -723 10629 -689 10663
rect -655 10629 -621 10663
rect -587 10629 -553 10663
rect -519 10629 -485 10663
rect -451 10629 -417 10663
rect -383 10629 -349 10663
rect -315 10629 -281 10663
rect -247 10629 -213 10663
rect -179 10629 -145 10663
rect -111 10629 -77 10663
rect -43 10629 -9 10663
rect 25 10629 59 10663
rect 93 10629 127 10663
rect 161 10629 195 10663
rect 229 10629 263 10663
rect 297 10629 331 10663
rect 365 10629 457 10663
rect -1353 10551 -1319 10629
rect -1193 10527 -1146 10561
rect -1110 10527 -1076 10561
rect -1040 10527 -993 10561
rect 97 10527 144 10561
rect 180 10527 214 10561
rect 250 10527 297 10561
rect 423 10551 457 10629
rect -1353 10483 -1319 10517
rect -1353 10415 -1319 10449
rect -1353 10347 -1319 10381
rect -1353 10279 -1319 10313
rect -1239 10465 -1205 10484
rect -1239 10397 -1205 10399
rect -1239 10361 -1205 10363
rect -1239 10276 -1205 10295
rect -981 10465 -947 10484
rect -981 10397 -947 10399
rect -981 10361 -947 10363
rect -981 10276 -947 10295
rect -723 10465 -689 10484
rect -723 10397 -689 10399
rect -723 10361 -689 10363
rect -723 10276 -689 10295
rect -465 10465 -431 10484
rect -465 10397 -431 10399
rect -465 10361 -431 10363
rect -465 10276 -431 10295
rect -207 10465 -173 10484
rect -207 10397 -173 10399
rect -207 10361 -173 10363
rect -207 10276 -173 10295
rect 51 10465 85 10484
rect 51 10397 85 10399
rect 51 10361 85 10363
rect 51 10276 85 10295
rect 309 10465 343 10484
rect 309 10397 343 10399
rect 309 10361 343 10363
rect 309 10276 343 10295
rect 423 10483 457 10517
rect 423 10415 457 10449
rect 423 10347 457 10381
rect 423 10279 457 10313
rect -1353 10211 -1319 10245
rect -1193 10199 -1146 10233
rect -1110 10199 -1076 10233
rect -1040 10199 -993 10233
rect -935 10199 -888 10233
rect -852 10199 -818 10233
rect -782 10199 -735 10233
rect -677 10199 -630 10233
rect -594 10199 -560 10233
rect -524 10199 -477 10233
rect -419 10199 -372 10233
rect -336 10199 -302 10233
rect -266 10199 -219 10233
rect -161 10199 -114 10233
rect -78 10199 -44 10233
rect -8 10199 39 10233
rect 97 10199 144 10233
rect 180 10199 214 10233
rect 250 10199 297 10233
rect 423 10211 457 10245
rect -1353 10143 -1319 10177
rect 423 10143 457 10177
rect -1353 10075 -1319 10109
rect -1193 10091 -1146 10125
rect -1110 10091 -1076 10125
rect -1040 10091 -993 10125
rect -935 10091 -888 10125
rect -852 10091 -818 10125
rect -782 10091 -735 10125
rect -677 10091 -630 10125
rect -594 10091 -560 10125
rect -524 10091 -477 10125
rect -419 10091 -372 10125
rect -336 10091 -302 10125
rect -266 10091 -219 10125
rect -161 10091 -114 10125
rect -78 10091 -44 10125
rect -8 10091 39 10125
rect 97 10091 144 10125
rect 180 10091 214 10125
rect 250 10091 297 10125
rect 423 10075 457 10109
rect -1353 10007 -1319 10041
rect -1353 9939 -1319 9973
rect -1353 9871 -1319 9905
rect -1239 10029 -1205 10048
rect -1239 9961 -1205 9963
rect -1239 9925 -1205 9927
rect -1239 9840 -1205 9859
rect -981 10029 -947 10048
rect -981 9961 -947 9963
rect -981 9925 -947 9927
rect -981 9840 -947 9859
rect -723 10029 -689 10048
rect -723 9961 -689 9963
rect -723 9925 -689 9927
rect -723 9840 -689 9859
rect -465 10029 -431 10048
rect -465 9961 -431 9963
rect -465 9925 -431 9927
rect -465 9840 -431 9859
rect -207 10029 -173 10048
rect -207 9961 -173 9963
rect -207 9925 -173 9927
rect -207 9840 -173 9859
rect 51 10029 85 10048
rect 51 9961 85 9963
rect 51 9925 85 9927
rect 51 9840 85 9859
rect 309 10029 343 10048
rect 309 9961 343 9963
rect 309 9925 343 9927
rect 309 9840 343 9859
rect 423 10007 457 10041
rect 423 9939 457 9973
rect 423 9871 457 9905
rect -1353 9803 -1319 9837
rect 423 9803 457 9837
rect -1353 9735 -1319 9769
rect -1193 9763 -1146 9797
rect -1110 9763 -1076 9797
rect -1040 9763 -993 9797
rect 97 9763 144 9797
rect 180 9763 214 9797
rect 250 9763 297 9797
rect -1353 9667 -1319 9701
rect 423 9735 457 9769
rect -1193 9655 -1146 9689
rect -1110 9655 -1076 9689
rect -1040 9655 -993 9689
rect 97 9655 144 9689
rect 180 9655 214 9689
rect 250 9655 297 9689
rect 423 9667 457 9701
rect -1353 9599 -1319 9633
rect -1353 9531 -1319 9565
rect -1353 9463 -1319 9497
rect -1353 9395 -1319 9429
rect -1239 9593 -1205 9612
rect -1239 9525 -1205 9527
rect -1239 9489 -1205 9491
rect -1239 9404 -1205 9423
rect -981 9593 -947 9612
rect -981 9525 -947 9527
rect -981 9489 -947 9491
rect -981 9404 -947 9423
rect -723 9593 -689 9612
rect -723 9525 -689 9527
rect -723 9489 -689 9491
rect -723 9404 -689 9423
rect -465 9593 -431 9612
rect -465 9525 -431 9527
rect -465 9489 -431 9491
rect -465 9404 -431 9423
rect -207 9593 -173 9612
rect -207 9525 -173 9527
rect -207 9489 -173 9491
rect -207 9404 -173 9423
rect 51 9593 85 9612
rect 51 9525 85 9527
rect 51 9489 85 9491
rect 51 9404 85 9423
rect 309 9593 343 9612
rect 309 9525 343 9527
rect 309 9489 343 9491
rect 309 9404 343 9423
rect 423 9599 457 9633
rect 423 9531 457 9565
rect 423 9463 457 9497
rect 423 9395 457 9429
rect -1353 9327 -1319 9361
rect -1193 9327 -1146 9361
rect -1110 9327 -1076 9361
rect -1040 9327 -993 9361
rect -935 9327 -888 9361
rect -852 9327 -818 9361
rect -782 9327 -735 9361
rect -677 9327 -630 9361
rect -594 9327 -560 9361
rect -524 9327 -477 9361
rect -419 9327 -372 9361
rect -336 9327 -302 9361
rect -266 9327 -219 9361
rect -161 9327 -114 9361
rect -78 9327 -44 9361
rect -8 9327 39 9361
rect 97 9327 144 9361
rect 180 9327 214 9361
rect 250 9327 297 9361
rect 423 9327 457 9361
rect -1353 9259 -1319 9293
rect 423 9259 457 9293
rect -1353 9191 -1319 9225
rect -1193 9219 -1146 9253
rect -1110 9219 -1076 9253
rect -1040 9219 -993 9253
rect -935 9219 -888 9253
rect -852 9219 -818 9253
rect -782 9219 -735 9253
rect -677 9219 -630 9253
rect -594 9219 -560 9253
rect -524 9219 -477 9253
rect -419 9219 -372 9253
rect -336 9219 -302 9253
rect -266 9219 -219 9253
rect -161 9219 -114 9253
rect -78 9219 -44 9253
rect -8 9219 39 9253
rect 97 9219 144 9253
rect 180 9219 214 9253
rect 250 9219 297 9253
rect 423 9191 457 9225
rect -1353 9123 -1319 9157
rect -1353 9055 -1319 9089
rect -1353 8987 -1319 9021
rect -1239 9157 -1205 9176
rect -1239 9089 -1205 9091
rect -1239 9053 -1205 9055
rect -1239 8968 -1205 8987
rect -981 9157 -947 9176
rect -981 9089 -947 9091
rect -981 9053 -947 9055
rect -981 8968 -947 8987
rect -723 9157 -689 9176
rect -723 9089 -689 9091
rect -723 9053 -689 9055
rect -723 8968 -689 8987
rect -465 9157 -431 9176
rect -465 9089 -431 9091
rect -465 9053 -431 9055
rect -465 8968 -431 8987
rect -207 9157 -173 9176
rect -207 9089 -173 9091
rect -207 9053 -173 9055
rect -207 8968 -173 8987
rect 51 9157 85 9176
rect 51 9089 85 9091
rect 51 9053 85 9055
rect 51 8968 85 8987
rect 309 9157 343 9176
rect 309 9089 343 9091
rect 309 9053 343 9055
rect 309 8968 343 8987
rect 423 9123 457 9157
rect 423 9055 457 9089
rect 423 8987 457 9021
rect -1353 8919 -1319 8953
rect -1193 8891 -1146 8925
rect -1110 8891 -1076 8925
rect -1040 8891 -993 8925
rect 97 8891 144 8925
rect 180 8891 214 8925
rect 250 8891 297 8925
rect 423 8919 457 8953
rect -1353 8823 -1319 8885
rect 423 8823 457 8885
rect -1353 8789 -1233 8823
rect -1199 8789 -1165 8823
rect -1131 8789 -1097 8823
rect -1063 8789 -1029 8823
rect -995 8789 -961 8823
rect -927 8789 -893 8823
rect -859 8789 -825 8823
rect -791 8789 -757 8823
rect -723 8789 -689 8823
rect -655 8789 -621 8823
rect -587 8789 -553 8823
rect -519 8789 -485 8823
rect -451 8789 -417 8823
rect -383 8789 -349 8823
rect -315 8789 -281 8823
rect -247 8789 -213 8823
rect -179 8789 -145 8823
rect -111 8789 -77 8823
rect -43 8789 -9 8823
rect 25 8789 59 8823
rect 93 8789 127 8823
rect 161 8789 195 8823
rect 229 8789 263 8823
rect 297 8789 331 8823
rect 365 8789 457 8823
rect 2969 10635 3003 10669
rect 2969 10567 3003 10601
rect 2969 10499 3003 10533
rect 3083 10684 3117 10703
rect 3083 10616 3117 10618
rect 3083 10580 3117 10582
rect 3083 10495 3117 10514
rect 3341 10684 3375 10703
rect 3341 10616 3375 10618
rect 3341 10580 3375 10582
rect 3341 10495 3375 10514
rect 3599 10684 3633 10703
rect 3599 10616 3633 10618
rect 3599 10580 3633 10582
rect 3599 10495 3633 10514
rect 3857 10684 3891 10703
rect 3857 10616 3891 10618
rect 3857 10580 3891 10582
rect 3857 10495 3891 10514
rect 4115 10684 4149 10703
rect 4115 10616 4149 10618
rect 4115 10580 4149 10582
rect 4115 10495 4149 10514
rect 4373 10684 4407 10703
rect 4373 10616 4407 10618
rect 4373 10580 4407 10582
rect 4373 10495 4407 10514
rect 4631 10684 4665 10703
rect 4631 10616 4665 10618
rect 4631 10580 4665 10582
rect 4631 10495 4665 10514
rect 4889 10684 4923 10703
rect 4889 10616 4923 10618
rect 4889 10580 4923 10582
rect 4889 10495 4923 10514
rect 5147 10684 5181 10703
rect 5147 10616 5181 10618
rect 5147 10580 5181 10582
rect 5147 10495 5181 10514
rect 5262 10635 5296 10669
rect 5262 10567 5296 10601
rect 5262 10499 5296 10533
rect 2969 10431 3003 10465
rect 3129 10427 3176 10461
rect 3212 10427 3246 10461
rect 3282 10427 3329 10461
rect 3903 10427 3950 10461
rect 3986 10427 4020 10461
rect 4056 10427 4103 10461
rect 4161 10427 4208 10461
rect 4244 10427 4278 10461
rect 4314 10427 4361 10461
rect 4935 10424 4982 10458
rect 5018 10424 5052 10458
rect 5088 10424 5135 10458
rect 5262 10431 5296 10465
rect 2969 10363 3003 10397
rect 5262 10363 5296 10397
rect 2969 10295 3003 10329
rect 3129 10319 3176 10353
rect 3212 10319 3246 10353
rect 3282 10319 3329 10353
rect 3903 10319 3950 10353
rect 3986 10319 4020 10353
rect 4056 10319 4103 10353
rect 4161 10319 4208 10353
rect 4244 10319 4278 10353
rect 4314 10319 4361 10353
rect 4935 10319 4982 10353
rect 5018 10319 5052 10353
rect 5088 10319 5135 10353
rect 5262 10295 5296 10329
rect 2969 10227 3003 10261
rect 2969 10159 3003 10193
rect 2969 10091 3003 10125
rect 3083 10266 3117 10285
rect 3083 10198 3117 10200
rect 3083 10162 3117 10164
rect 3083 10077 3117 10096
rect 3341 10266 3375 10285
rect 3341 10198 3375 10200
rect 3341 10162 3375 10164
rect 3341 10077 3375 10096
rect 3599 10266 3633 10285
rect 3599 10198 3633 10200
rect 3599 10162 3633 10164
rect 3599 10077 3633 10096
rect 3857 10266 3891 10285
rect 3857 10198 3891 10200
rect 3857 10162 3891 10164
rect 3857 10077 3891 10096
rect 4115 10266 4149 10285
rect 4115 10198 4149 10200
rect 4115 10162 4149 10164
rect 4115 10077 4149 10096
rect 4373 10266 4407 10285
rect 4373 10198 4407 10200
rect 4373 10162 4407 10164
rect 4373 10077 4407 10096
rect 4631 10266 4665 10285
rect 4631 10198 4665 10200
rect 4631 10162 4665 10164
rect 4631 10077 4665 10096
rect 4889 10266 4923 10285
rect 4889 10198 4923 10200
rect 4889 10162 4923 10164
rect 4889 10077 4923 10096
rect 5147 10266 5181 10285
rect 5147 10198 5181 10200
rect 5147 10162 5181 10164
rect 5147 10077 5181 10096
rect 5262 10227 5296 10261
rect 5262 10159 5296 10193
rect 5262 10091 5296 10125
rect 2969 10023 3003 10057
rect 3129 10009 3176 10043
rect 3212 10009 3246 10043
rect 3282 10009 3329 10043
rect 3387 10009 3434 10043
rect 3470 10009 3504 10043
rect 3540 10009 3587 10043
rect 3645 10009 3692 10043
rect 3728 10009 3762 10043
rect 3798 10009 3845 10043
rect 4419 10009 4466 10043
rect 4502 10009 4536 10043
rect 4572 10009 4619 10043
rect 4677 10009 4724 10043
rect 4760 10009 4794 10043
rect 4830 10009 4877 10043
rect 4935 10009 4982 10043
rect 5018 10009 5052 10043
rect 5088 10009 5135 10043
rect 5262 10023 5296 10057
rect 2969 9955 3003 9989
rect 5262 9955 5296 9989
rect 2969 9887 3003 9921
rect 3129 9901 3176 9935
rect 3212 9901 3246 9935
rect 3282 9901 3329 9935
rect 3387 9901 3434 9935
rect 3470 9901 3504 9935
rect 3540 9901 3587 9935
rect 3645 9901 3692 9935
rect 3728 9901 3762 9935
rect 3798 9901 3845 9935
rect 4419 9901 4466 9935
rect 4502 9901 4536 9935
rect 4572 9901 4619 9935
rect 4677 9901 4724 9935
rect 4760 9901 4794 9935
rect 4830 9901 4877 9935
rect 4935 9901 4982 9935
rect 5018 9901 5052 9935
rect 5088 9901 5135 9935
rect 5262 9887 5296 9921
rect 2969 9819 3003 9853
rect 2969 9751 3003 9785
rect 2969 9683 3003 9717
rect 3083 9848 3117 9867
rect 3083 9780 3117 9782
rect 3083 9744 3117 9746
rect 3083 9659 3117 9678
rect 3341 9848 3375 9867
rect 3341 9780 3375 9782
rect 3341 9744 3375 9746
rect 3341 9659 3375 9678
rect 3599 9848 3633 9867
rect 3599 9780 3633 9782
rect 3599 9744 3633 9746
rect 3599 9659 3633 9678
rect 3857 9848 3891 9867
rect 3857 9780 3891 9782
rect 3857 9744 3891 9746
rect 3857 9659 3891 9678
rect 4115 9848 4149 9867
rect 4115 9780 4149 9782
rect 4115 9744 4149 9746
rect 4115 9659 4149 9678
rect 4373 9848 4407 9867
rect 4373 9780 4407 9782
rect 4373 9744 4407 9746
rect 4373 9659 4407 9678
rect 4631 9848 4665 9867
rect 4631 9780 4665 9782
rect 4631 9744 4665 9746
rect 4631 9659 4665 9678
rect 4889 9848 4923 9867
rect 4889 9780 4923 9782
rect 4889 9744 4923 9746
rect 4889 9659 4923 9678
rect 5147 9848 5181 9867
rect 5147 9780 5181 9782
rect 5147 9744 5181 9746
rect 5147 9659 5181 9678
rect 5262 9819 5296 9853
rect 5262 9751 5296 9785
rect 5262 9683 5296 9717
rect 2969 9615 3003 9649
rect 3129 9591 3176 9625
rect 3212 9591 3246 9625
rect 3282 9591 3329 9625
rect 3903 9591 3950 9625
rect 3986 9591 4020 9625
rect 4056 9591 4103 9625
rect 4161 9591 4208 9625
rect 4244 9591 4278 9625
rect 4314 9591 4361 9625
rect 4935 9588 4982 9622
rect 5018 9588 5052 9622
rect 5088 9588 5135 9622
rect 5262 9615 5296 9649
rect 2969 9547 3003 9581
rect 5262 9547 5296 9581
rect 2969 9479 3003 9513
rect 3129 9483 3176 9517
rect 3212 9483 3246 9517
rect 3282 9483 3329 9517
rect 3903 9483 3950 9517
rect 3986 9483 4020 9517
rect 4056 9483 4103 9517
rect 4161 9483 4208 9517
rect 4244 9483 4278 9517
rect 4314 9483 4361 9517
rect 4935 9483 4982 9517
rect 5018 9483 5052 9517
rect 5088 9483 5135 9517
rect 5262 9479 5296 9513
rect 2969 9411 3003 9445
rect 2969 9343 3003 9377
rect 2969 9275 3003 9309
rect 3083 9430 3117 9449
rect 3083 9362 3117 9364
rect 3083 9326 3117 9328
rect 3083 9241 3117 9260
rect 3341 9430 3375 9449
rect 3341 9362 3375 9364
rect 3341 9326 3375 9328
rect 3341 9241 3375 9260
rect 3599 9430 3633 9449
rect 3599 9362 3633 9364
rect 3599 9326 3633 9328
rect 3599 9241 3633 9260
rect 3857 9430 3891 9449
rect 3857 9362 3891 9364
rect 3857 9326 3891 9328
rect 3857 9241 3891 9260
rect 4115 9430 4149 9449
rect 4115 9362 4149 9364
rect 4115 9326 4149 9328
rect 4115 9241 4149 9260
rect 4373 9430 4407 9449
rect 4373 9362 4407 9364
rect 4373 9326 4407 9328
rect 4373 9241 4407 9260
rect 4631 9430 4665 9449
rect 4631 9362 4665 9364
rect 4631 9326 4665 9328
rect 4631 9241 4665 9260
rect 4889 9430 4923 9449
rect 4889 9362 4923 9364
rect 4889 9326 4923 9328
rect 4889 9241 4923 9260
rect 5147 9430 5181 9449
rect 5147 9362 5181 9364
rect 5147 9326 5181 9328
rect 5147 9241 5181 9260
rect 5262 9411 5296 9445
rect 5262 9343 5296 9377
rect 5262 9275 5296 9309
rect 2969 9207 3003 9241
rect 5262 9207 5296 9241
rect 3129 9173 3176 9207
rect 3212 9173 3246 9207
rect 3282 9173 3329 9207
rect 3387 9173 3434 9207
rect 3470 9173 3504 9207
rect 3540 9173 3587 9207
rect 3645 9173 3692 9207
rect 3728 9173 3762 9207
rect 3798 9173 3845 9207
rect 4419 9173 4466 9207
rect 4502 9173 4536 9207
rect 4572 9173 4619 9207
rect 4677 9173 4724 9207
rect 4760 9173 4794 9207
rect 4830 9173 4877 9207
rect 2969 9139 3003 9173
rect 4935 9170 4982 9204
rect 5018 9170 5052 9204
rect 5088 9170 5135 9204
rect 2969 9071 3003 9105
rect 5262 9139 5296 9173
rect 3129 9061 3176 9095
rect 3212 9061 3246 9095
rect 3282 9061 3329 9095
rect 3387 9061 3434 9095
rect 3470 9061 3504 9095
rect 3540 9061 3587 9095
rect 3645 9061 3692 9095
rect 3728 9061 3762 9095
rect 3798 9061 3845 9095
rect 4419 9061 4466 9095
rect 4502 9061 4536 9095
rect 4572 9061 4619 9095
rect 4677 9061 4724 9095
rect 4760 9061 4794 9095
rect 4830 9061 4877 9095
rect 4935 9061 4982 9095
rect 5018 9061 5052 9095
rect 5088 9061 5135 9095
rect 5262 9071 5296 9105
rect 2969 9003 3003 9037
rect 2969 8935 3003 8969
rect 2969 8867 3003 8901
rect 2969 8799 3003 8833
rect 3083 9008 3117 9027
rect 3083 8940 3117 8942
rect 3083 8904 3117 8906
rect 3083 8819 3117 8838
rect 3341 9008 3375 9027
rect 3341 8940 3375 8942
rect 3341 8904 3375 8906
rect 3341 8819 3375 8838
rect 3599 9008 3633 9027
rect 3599 8940 3633 8942
rect 3599 8904 3633 8906
rect 3599 8819 3633 8838
rect 3857 9008 3891 9027
rect 3857 8940 3891 8942
rect 3857 8904 3891 8906
rect 3857 8819 3891 8838
rect 4115 9008 4149 9027
rect 4115 8940 4149 8942
rect 4115 8904 4149 8906
rect 4115 8819 4149 8838
rect 4373 9008 4407 9027
rect 4373 8940 4407 8942
rect 4373 8904 4407 8906
rect 4373 8819 4407 8838
rect 4631 9008 4665 9027
rect 4631 8940 4665 8942
rect 4631 8904 4665 8906
rect 4631 8819 4665 8838
rect 4889 9008 4923 9027
rect 4889 8940 4923 8942
rect 4889 8904 4923 8906
rect 4889 8819 4923 8838
rect 5147 9008 5181 9027
rect 5147 8940 5181 8942
rect 5147 8904 5181 8906
rect 5147 8819 5181 8838
rect 5262 9003 5296 9037
rect 5262 8935 5296 8969
rect 5262 8867 5296 8901
rect 5262 8799 5296 8833
rect 2969 8731 3003 8765
rect 3129 8751 3176 8785
rect 3212 8751 3246 8785
rect 3282 8751 3329 8785
rect 3903 8751 3950 8785
rect 3986 8751 4020 8785
rect 4056 8751 4103 8785
rect 4161 8751 4208 8785
rect 4244 8751 4278 8785
rect 4314 8751 4361 8785
rect 4935 8748 4982 8782
rect 5018 8748 5052 8782
rect 5088 8748 5135 8782
rect 2969 8663 3003 8697
rect 5262 8731 5296 8765
rect 3129 8639 3176 8673
rect 3212 8639 3246 8673
rect 3282 8639 3329 8673
rect 3903 8639 3950 8673
rect 3986 8639 4020 8673
rect 4056 8639 4103 8673
rect 4161 8639 4208 8673
rect 4244 8639 4278 8673
rect 4314 8639 4361 8673
rect 4935 8639 4982 8673
rect 5018 8639 5052 8673
rect 5088 8639 5135 8673
rect 5262 8663 5296 8697
rect 2969 8595 3003 8629
rect 2969 8527 3003 8561
rect 2969 8459 3003 8493
rect 2969 8391 3003 8425
rect 3083 8586 3117 8605
rect 3083 8518 3117 8520
rect 3083 8482 3117 8484
rect 3083 8397 3117 8416
rect 3341 8586 3375 8605
rect 3341 8518 3375 8520
rect 3341 8482 3375 8484
rect 3341 8397 3375 8416
rect 3599 8586 3633 8605
rect 3599 8518 3633 8520
rect 3599 8482 3633 8484
rect 3599 8397 3633 8416
rect 3857 8586 3891 8605
rect 3857 8518 3891 8520
rect 3857 8482 3891 8484
rect 3857 8397 3891 8416
rect 4115 8586 4149 8605
rect 4115 8518 4149 8520
rect 4115 8482 4149 8484
rect 4115 8397 4149 8416
rect 4373 8586 4407 8605
rect 4373 8518 4407 8520
rect 4373 8482 4407 8484
rect 4373 8397 4407 8416
rect 4631 8586 4665 8605
rect 4631 8518 4665 8520
rect 4631 8482 4665 8484
rect 4631 8397 4665 8416
rect 4889 8586 4923 8605
rect 4889 8518 4923 8520
rect 4889 8482 4923 8484
rect 4889 8397 4923 8416
rect 5147 8586 5181 8605
rect 5147 8518 5181 8520
rect 5147 8482 5181 8484
rect 5147 8397 5181 8416
rect 5262 8595 5296 8629
rect 5262 8527 5296 8561
rect 5262 8459 5296 8493
rect 5262 8391 5296 8425
rect 3129 8329 3176 8363
rect 3212 8329 3246 8363
rect 3282 8329 3329 8363
rect 3387 8329 3434 8363
rect 3470 8329 3504 8363
rect 3540 8329 3587 8363
rect 3645 8329 3692 8363
rect 3728 8329 3762 8363
rect 3798 8329 3845 8363
rect 4419 8329 4466 8363
rect 4502 8329 4536 8363
rect 4572 8329 4619 8363
rect 4677 8329 4724 8363
rect 4760 8329 4794 8363
rect 4830 8329 4877 8363
rect 4935 8329 4982 8363
rect 5018 8329 5052 8363
rect 5088 8329 5135 8363
rect 2969 8268 3003 8329
rect 5262 8268 5296 8357
rect 2969 8234 3089 8268
rect 3123 8234 3157 8268
rect 3191 8234 3225 8268
rect 3259 8234 3293 8268
rect 3327 8234 3361 8268
rect 3395 8234 3429 8268
rect 3463 8234 3497 8268
rect 3531 8234 3565 8268
rect 3599 8234 3633 8268
rect 3667 8234 3701 8268
rect 3735 8234 3769 8268
rect 3803 8234 3837 8268
rect 3871 8234 3905 8268
rect 3939 8234 3973 8268
rect 4007 8234 4041 8268
rect 4075 8234 4109 8268
rect 4143 8234 4177 8268
rect 4211 8234 4245 8268
rect 4279 8234 4313 8268
rect 4347 8234 4381 8268
rect 4415 8234 4449 8268
rect 4483 8234 4517 8268
rect 4551 8234 4585 8268
rect 4619 8234 4653 8268
rect 4687 8234 4721 8268
rect 4755 8234 4789 8268
rect 4823 8234 4857 8268
rect 4891 8234 4925 8268
rect 4959 8234 4993 8268
rect 5027 8234 5061 8268
rect 5095 8234 5129 8268
rect 5163 8234 5296 8268
rect 6895 10869 6929 10947
rect 7055 10845 7102 10879
rect 7138 10845 7172 10879
rect 7208 10845 7255 10879
rect 8345 10845 8392 10879
rect 8428 10845 8462 10879
rect 8498 10845 8545 10879
rect 8671 10869 8705 10947
rect 6895 10801 6929 10835
rect 6895 10733 6929 10767
rect 6895 10665 6929 10699
rect 6895 10597 6929 10631
rect 7009 10783 7043 10802
rect 7009 10715 7043 10717
rect 7009 10679 7043 10681
rect 7009 10594 7043 10613
rect 7267 10783 7301 10802
rect 7267 10715 7301 10717
rect 7267 10679 7301 10681
rect 7267 10594 7301 10613
rect 7525 10783 7559 10802
rect 7525 10715 7559 10717
rect 7525 10679 7559 10681
rect 7525 10594 7559 10613
rect 7783 10783 7817 10802
rect 7783 10715 7817 10717
rect 7783 10679 7817 10681
rect 7783 10594 7817 10613
rect 8041 10783 8075 10802
rect 8041 10715 8075 10717
rect 8041 10679 8075 10681
rect 8041 10594 8075 10613
rect 8299 10783 8333 10802
rect 8299 10715 8333 10717
rect 8299 10679 8333 10681
rect 8299 10594 8333 10613
rect 8557 10783 8591 10802
rect 8557 10715 8591 10717
rect 8557 10679 8591 10681
rect 8557 10594 8591 10613
rect 8671 10801 8705 10835
rect 8671 10733 8705 10767
rect 8671 10665 8705 10699
rect 8671 10597 8705 10631
rect 6895 10529 6929 10563
rect 7055 10517 7102 10551
rect 7138 10517 7172 10551
rect 7208 10517 7255 10551
rect 7313 10517 7360 10551
rect 7396 10517 7430 10551
rect 7466 10517 7513 10551
rect 7571 10517 7618 10551
rect 7654 10517 7688 10551
rect 7724 10517 7771 10551
rect 7829 10517 7876 10551
rect 7912 10517 7946 10551
rect 7982 10517 8029 10551
rect 8087 10517 8134 10551
rect 8170 10517 8204 10551
rect 8240 10517 8287 10551
rect 8345 10517 8392 10551
rect 8428 10517 8462 10551
rect 8498 10517 8545 10551
rect 8671 10529 8705 10563
rect 6895 10461 6929 10495
rect 8671 10461 8705 10495
rect 6895 10393 6929 10427
rect 7055 10409 7102 10443
rect 7138 10409 7172 10443
rect 7208 10409 7255 10443
rect 7313 10409 7360 10443
rect 7396 10409 7430 10443
rect 7466 10409 7513 10443
rect 7571 10409 7618 10443
rect 7654 10409 7688 10443
rect 7724 10409 7771 10443
rect 7829 10409 7876 10443
rect 7912 10409 7946 10443
rect 7982 10409 8029 10443
rect 8087 10409 8134 10443
rect 8170 10409 8204 10443
rect 8240 10409 8287 10443
rect 8345 10409 8392 10443
rect 8428 10409 8462 10443
rect 8498 10409 8545 10443
rect 8671 10393 8705 10427
rect 6895 10325 6929 10359
rect 6895 10257 6929 10291
rect 6895 10189 6929 10223
rect 7009 10347 7043 10366
rect 7009 10279 7043 10281
rect 7009 10243 7043 10245
rect 7009 10158 7043 10177
rect 7267 10347 7301 10366
rect 7267 10279 7301 10281
rect 7267 10243 7301 10245
rect 7267 10158 7301 10177
rect 7525 10347 7559 10366
rect 7525 10279 7559 10281
rect 7525 10243 7559 10245
rect 7525 10158 7559 10177
rect 7783 10347 7817 10366
rect 7783 10279 7817 10281
rect 7783 10243 7817 10245
rect 7783 10158 7817 10177
rect 8041 10347 8075 10366
rect 8041 10279 8075 10281
rect 8041 10243 8075 10245
rect 8041 10158 8075 10177
rect 8299 10347 8333 10366
rect 8299 10279 8333 10281
rect 8299 10243 8333 10245
rect 8299 10158 8333 10177
rect 8557 10347 8591 10366
rect 8557 10279 8591 10281
rect 8557 10243 8591 10245
rect 8557 10158 8591 10177
rect 8671 10325 8705 10359
rect 8671 10257 8705 10291
rect 8671 10189 8705 10223
rect 6895 10121 6929 10155
rect 8671 10121 8705 10155
rect 6895 10053 6929 10087
rect 7055 10081 7102 10115
rect 7138 10081 7172 10115
rect 7208 10081 7255 10115
rect 8345 10081 8392 10115
rect 8428 10081 8462 10115
rect 8498 10081 8545 10115
rect 6895 9985 6929 10019
rect 8671 10053 8705 10087
rect 7055 9973 7102 10007
rect 7138 9973 7172 10007
rect 7208 9973 7255 10007
rect 8345 9973 8392 10007
rect 8428 9973 8462 10007
rect 8498 9973 8545 10007
rect 8671 9985 8705 10019
rect 6895 9917 6929 9951
rect 6895 9849 6929 9883
rect 6895 9781 6929 9815
rect 6895 9713 6929 9747
rect 7009 9911 7043 9930
rect 7009 9843 7043 9845
rect 7009 9807 7043 9809
rect 7009 9722 7043 9741
rect 7267 9911 7301 9930
rect 7267 9843 7301 9845
rect 7267 9807 7301 9809
rect 7267 9722 7301 9741
rect 7525 9911 7559 9930
rect 7525 9843 7559 9845
rect 7525 9807 7559 9809
rect 7525 9722 7559 9741
rect 7783 9911 7817 9930
rect 7783 9843 7817 9845
rect 7783 9807 7817 9809
rect 7783 9722 7817 9741
rect 8041 9911 8075 9930
rect 8041 9843 8075 9845
rect 8041 9807 8075 9809
rect 8041 9722 8075 9741
rect 8299 9911 8333 9930
rect 8299 9843 8333 9845
rect 8299 9807 8333 9809
rect 8299 9722 8333 9741
rect 8557 9911 8591 9930
rect 8557 9843 8591 9845
rect 8557 9807 8591 9809
rect 8557 9722 8591 9741
rect 8671 9917 8705 9951
rect 8671 9849 8705 9883
rect 8671 9781 8705 9815
rect 8671 9713 8705 9747
rect 6895 9645 6929 9679
rect 7055 9645 7102 9679
rect 7138 9645 7172 9679
rect 7208 9645 7255 9679
rect 7313 9645 7360 9679
rect 7396 9645 7430 9679
rect 7466 9645 7513 9679
rect 7571 9645 7618 9679
rect 7654 9645 7688 9679
rect 7724 9645 7771 9679
rect 7829 9645 7876 9679
rect 7912 9645 7946 9679
rect 7982 9645 8029 9679
rect 8087 9645 8134 9679
rect 8170 9645 8204 9679
rect 8240 9645 8287 9679
rect 8345 9645 8392 9679
rect 8428 9645 8462 9679
rect 8498 9645 8545 9679
rect 8671 9645 8705 9679
rect 6895 9577 6929 9611
rect 8671 9577 8705 9611
rect 6895 9509 6929 9543
rect 7055 9537 7102 9571
rect 7138 9537 7172 9571
rect 7208 9537 7255 9571
rect 7313 9537 7360 9571
rect 7396 9537 7430 9571
rect 7466 9537 7513 9571
rect 7571 9537 7618 9571
rect 7654 9537 7688 9571
rect 7724 9537 7771 9571
rect 7829 9537 7876 9571
rect 7912 9537 7946 9571
rect 7982 9537 8029 9571
rect 8087 9537 8134 9571
rect 8170 9537 8204 9571
rect 8240 9537 8287 9571
rect 8345 9537 8392 9571
rect 8428 9537 8462 9571
rect 8498 9537 8545 9571
rect 8671 9509 8705 9543
rect 6895 9441 6929 9475
rect 6895 9373 6929 9407
rect 6895 9305 6929 9339
rect 7009 9475 7043 9494
rect 7009 9407 7043 9409
rect 7009 9371 7043 9373
rect 7009 9286 7043 9305
rect 7267 9475 7301 9494
rect 7267 9407 7301 9409
rect 7267 9371 7301 9373
rect 7267 9286 7301 9305
rect 7525 9475 7559 9494
rect 7525 9407 7559 9409
rect 7525 9371 7559 9373
rect 7525 9286 7559 9305
rect 7783 9475 7817 9494
rect 7783 9407 7817 9409
rect 7783 9371 7817 9373
rect 7783 9286 7817 9305
rect 8041 9475 8075 9494
rect 8041 9407 8075 9409
rect 8041 9371 8075 9373
rect 8041 9286 8075 9305
rect 8299 9475 8333 9494
rect 8299 9407 8333 9409
rect 8299 9371 8333 9373
rect 8299 9286 8333 9305
rect 8557 9475 8591 9494
rect 8557 9407 8591 9409
rect 8557 9371 8591 9373
rect 8557 9286 8591 9305
rect 8671 9441 8705 9475
rect 8671 9373 8705 9407
rect 8671 9305 8705 9339
rect 6895 9237 6929 9271
rect 7055 9209 7102 9243
rect 7138 9209 7172 9243
rect 7208 9209 7255 9243
rect 8345 9209 8392 9243
rect 8428 9209 8462 9243
rect 8498 9209 8545 9243
rect 8671 9237 8705 9271
rect 6895 9169 6929 9203
rect 8671 9169 8705 9203
rect 6895 9101 6929 9135
rect 7055 9101 7102 9135
rect 7138 9101 7172 9135
rect 7208 9101 7255 9135
rect 8345 9101 8392 9135
rect 8428 9101 8462 9135
rect 8498 9101 8545 9135
rect 8671 9101 8705 9135
rect 6895 9033 6929 9067
rect 6895 8965 6929 8999
rect 6895 8897 6929 8931
rect 6895 8829 6929 8863
rect 7009 9039 7043 9058
rect 7009 8971 7043 8973
rect 7009 8935 7043 8937
rect 7009 8850 7043 8869
rect 7267 9039 7301 9058
rect 7267 8971 7301 8973
rect 7267 8935 7301 8937
rect 7267 8850 7301 8869
rect 7525 9039 7559 9058
rect 7525 8971 7559 8973
rect 7525 8935 7559 8937
rect 7525 8850 7559 8869
rect 7783 9039 7817 9058
rect 7783 8971 7817 8973
rect 7783 8935 7817 8937
rect 7783 8850 7817 8869
rect 8041 9039 8075 9058
rect 8041 8971 8075 8973
rect 8041 8935 8075 8937
rect 8041 8850 8075 8869
rect 8299 9039 8333 9058
rect 8299 8971 8333 8973
rect 8299 8935 8333 8937
rect 8299 8850 8333 8869
rect 8557 9039 8591 9058
rect 8557 8971 8591 8973
rect 8557 8935 8591 8937
rect 8557 8850 8591 8869
rect 8671 9033 8705 9067
rect 8671 8965 8705 8999
rect 8671 8897 8705 8931
rect 8671 8829 8705 8863
rect 6895 8761 6929 8795
rect 7055 8773 7102 8807
rect 7138 8773 7172 8807
rect 7208 8773 7255 8807
rect 7313 8773 7360 8807
rect 7396 8773 7430 8807
rect 7466 8773 7513 8807
rect 7571 8773 7618 8807
rect 7654 8773 7688 8807
rect 7724 8773 7771 8807
rect 7829 8773 7876 8807
rect 7912 8773 7946 8807
rect 7982 8773 8029 8807
rect 8087 8773 8134 8807
rect 8170 8773 8204 8807
rect 8240 8773 8287 8807
rect 8345 8773 8392 8807
rect 8428 8773 8462 8807
rect 8498 8773 8545 8807
rect 6895 8693 6929 8727
rect 8671 8761 8705 8795
rect 7055 8665 7102 8699
rect 7138 8665 7172 8699
rect 7208 8665 7255 8699
rect 7313 8665 7360 8699
rect 7396 8665 7430 8699
rect 7466 8665 7513 8699
rect 7571 8665 7618 8699
rect 7654 8665 7688 8699
rect 7724 8665 7771 8699
rect 7829 8665 7876 8699
rect 7912 8665 7946 8699
rect 7982 8665 8029 8699
rect 8087 8665 8134 8699
rect 8170 8665 8204 8699
rect 8240 8665 8287 8699
rect 8345 8665 8392 8699
rect 8428 8665 8462 8699
rect 8498 8665 8545 8699
rect 8671 8693 8705 8727
rect 6895 8625 6929 8659
rect 8671 8625 8705 8659
rect 6895 8557 6929 8591
rect 6895 8489 6929 8523
rect 6895 8421 6929 8455
rect 7009 8603 7043 8622
rect 7009 8535 7043 8537
rect 7009 8499 7043 8501
rect 7009 8414 7043 8433
rect 7267 8603 7301 8622
rect 7267 8535 7301 8537
rect 7267 8499 7301 8501
rect 7267 8414 7301 8433
rect 7525 8603 7559 8622
rect 7525 8535 7559 8537
rect 7525 8499 7559 8501
rect 7525 8414 7559 8433
rect 7783 8603 7817 8622
rect 7783 8535 7817 8537
rect 7783 8499 7817 8501
rect 7783 8414 7817 8433
rect 8041 8603 8075 8622
rect 8041 8535 8075 8537
rect 8041 8499 8075 8501
rect 8041 8414 8075 8433
rect 8299 8603 8333 8622
rect 8299 8535 8333 8537
rect 8299 8499 8333 8501
rect 8299 8414 8333 8433
rect 8557 8603 8591 8622
rect 8557 8535 8591 8537
rect 8557 8499 8591 8501
rect 8557 8414 8591 8433
rect 8671 8557 8705 8591
rect 8671 8489 8705 8523
rect 8671 8421 8705 8455
rect 6895 8353 6929 8387
rect 7055 8337 7102 8371
rect 7138 8337 7172 8371
rect 7208 8337 7255 8371
rect 8345 8337 8392 8371
rect 8428 8337 8462 8371
rect 8498 8337 8545 8371
rect 8671 8353 8705 8387
rect 6895 8285 6929 8319
rect 8671 8285 8705 8319
rect 6895 8217 6929 8251
rect 7055 8229 7102 8263
rect 7138 8229 7172 8263
rect 7208 8229 7255 8263
rect 7313 8229 7360 8263
rect 7396 8229 7430 8263
rect 7466 8229 7513 8263
rect 7571 8229 7618 8263
rect 7654 8229 7688 8263
rect 7724 8229 7771 8263
rect 7829 8229 7876 8263
rect 7912 8229 7946 8263
rect 7982 8229 8029 8263
rect 8087 8229 8134 8263
rect 8170 8229 8204 8263
rect 8240 8229 8287 8263
rect 8345 8229 8392 8263
rect 8428 8229 8462 8263
rect 8498 8229 8545 8263
rect 8671 8217 8705 8251
rect 6895 8149 6929 8183
rect -2322 8090 -2202 8124
rect -2168 8090 -2134 8124
rect -2100 8090 -2066 8124
rect -2032 8090 -1998 8124
rect -1964 8090 -1930 8124
rect -1896 8090 -1862 8124
rect -1828 8090 -1794 8124
rect -1760 8090 -1726 8124
rect -1692 8090 -1658 8124
rect -1624 8090 -1590 8124
rect -1556 8090 -1522 8124
rect -1488 8090 -1454 8124
rect -1420 8090 -1386 8124
rect -1352 8090 -1318 8124
rect -1284 8090 -1250 8124
rect -1216 8090 -1182 8124
rect -1148 8090 -1114 8124
rect -1080 8090 -1046 8124
rect -1012 8090 -978 8124
rect -944 8090 -910 8124
rect -876 8090 -842 8124
rect -808 8090 -774 8124
rect -740 8090 -706 8124
rect -672 8090 -638 8124
rect -604 8090 -570 8124
rect -536 8090 -502 8124
rect -468 8090 -434 8124
rect -400 8090 -366 8124
rect -332 8090 -298 8124
rect -264 8090 -230 8124
rect -196 8090 -162 8124
rect -128 8090 -94 8124
rect -60 8090 -26 8124
rect 8 8090 42 8124
rect 76 8090 110 8124
rect 144 8090 178 8124
rect 212 8090 246 8124
rect 280 8090 314 8124
rect 348 8090 382 8124
rect 416 8090 450 8124
rect 484 8090 518 8124
rect 552 8090 586 8124
rect 620 8090 654 8124
rect 688 8090 722 8124
rect 756 8090 790 8124
rect 824 8090 858 8124
rect 892 8090 926 8124
rect 960 8090 994 8124
rect 1028 8090 1062 8124
rect 1096 8090 1142 8124
rect 1176 8090 1210 8124
rect 1244 8090 1278 8124
rect 1312 8090 1346 8124
rect 1380 8090 1414 8124
rect 1448 8090 1552 8124
rect -2322 8002 -2288 8090
rect -2162 7988 -2115 8022
rect -2079 7988 -2045 8022
rect -2009 7988 -1962 8022
rect -1904 7988 -1857 8022
rect -1821 7988 -1787 8022
rect -1751 7988 -1704 8022
rect -1646 7988 -1599 8022
rect -1563 7988 -1529 8022
rect -1493 7988 -1446 8022
rect -1388 7988 -1341 8022
rect -1305 7988 -1271 8022
rect -1235 7988 -1188 8022
rect -1130 7988 -1083 8022
rect -1047 7988 -1013 8022
rect -977 7988 -930 8022
rect -872 7988 -825 8022
rect -789 7988 -755 8022
rect -719 7988 -672 8022
rect -614 7988 -567 8022
rect -531 7988 -497 8022
rect -461 7988 -414 8022
rect -356 7988 -309 8022
rect -273 7988 -239 8022
rect -203 7988 -156 8022
rect -98 7988 -51 8022
rect -15 7988 19 8022
rect 55 7988 102 8022
rect 160 7988 207 8022
rect 243 7988 277 8022
rect 313 7988 360 8022
rect 418 7988 465 8022
rect 501 7988 535 8022
rect 571 7988 618 8022
rect 676 7988 723 8022
rect 759 7988 793 8022
rect 829 7988 876 8022
rect 934 7988 981 8022
rect 1017 7988 1051 8022
rect 1087 7988 1134 8022
rect 1192 7988 1239 8022
rect 1275 7988 1309 8022
rect 1345 7988 1392 8022
rect 1518 8002 1552 8090
rect -2322 7934 -2288 7968
rect -2322 7866 -2288 7900
rect -2322 7798 -2288 7832
rect -2322 7730 -2288 7764
rect -2208 7935 -2174 7954
rect -2208 7867 -2174 7869
rect -2208 7831 -2174 7833
rect -2208 7746 -2174 7765
rect -1950 7935 -1916 7954
rect -1950 7867 -1916 7869
rect -1950 7831 -1916 7833
rect -1950 7746 -1916 7765
rect -1692 7935 -1658 7954
rect -1692 7867 -1658 7869
rect -1692 7831 -1658 7833
rect -1692 7746 -1658 7765
rect -1434 7935 -1400 7954
rect -1434 7867 -1400 7869
rect -1434 7831 -1400 7833
rect -1434 7746 -1400 7765
rect -1176 7935 -1142 7954
rect -1176 7867 -1142 7869
rect -1176 7831 -1142 7833
rect -1176 7746 -1142 7765
rect -918 7935 -884 7954
rect -918 7867 -884 7869
rect -918 7831 -884 7833
rect -918 7746 -884 7765
rect -660 7935 -626 7954
rect -660 7867 -626 7869
rect -660 7831 -626 7833
rect -660 7746 -626 7765
rect -402 7935 -368 7954
rect -402 7867 -368 7869
rect -402 7831 -368 7833
rect -402 7746 -368 7765
rect -144 7935 -110 7954
rect -144 7867 -110 7869
rect -144 7831 -110 7833
rect -144 7746 -110 7765
rect 114 7935 148 7954
rect 114 7867 148 7869
rect 114 7831 148 7833
rect 114 7746 148 7765
rect 372 7935 406 7954
rect 372 7867 406 7869
rect 372 7831 406 7833
rect 372 7746 406 7765
rect 630 7935 664 7954
rect 630 7867 664 7869
rect 630 7831 664 7833
rect 630 7746 664 7765
rect 888 7935 922 7954
rect 888 7867 922 7869
rect 888 7831 922 7833
rect 888 7746 922 7765
rect 1146 7935 1180 7954
rect 1146 7867 1180 7869
rect 1146 7831 1180 7833
rect 1146 7746 1180 7765
rect 1404 7935 1438 7954
rect 1404 7867 1438 7869
rect 1404 7831 1438 7833
rect 1404 7746 1438 7765
rect 1518 7934 1552 7968
rect 1518 7866 1552 7900
rect 1518 7798 1552 7832
rect 6895 8081 6929 8115
rect 6895 8013 6929 8047
rect 6895 7945 6929 7979
rect 7009 8167 7043 8186
rect 7009 8099 7043 8101
rect 7009 8063 7043 8065
rect 7009 7978 7043 7997
rect 7267 8167 7301 8186
rect 7267 8099 7301 8101
rect 7267 8063 7301 8065
rect 7267 7978 7301 7997
rect 7525 8167 7559 8186
rect 7525 8099 7559 8101
rect 7525 8063 7559 8065
rect 7525 7978 7559 7997
rect 7783 8167 7817 8186
rect 7783 8099 7817 8101
rect 7783 8063 7817 8065
rect 7783 7978 7817 7997
rect 8041 8167 8075 8186
rect 8041 8099 8075 8101
rect 8041 8063 8075 8065
rect 8041 7978 8075 7997
rect 8299 8167 8333 8186
rect 8299 8099 8333 8101
rect 8299 8063 8333 8065
rect 8299 7978 8333 7997
rect 8557 8167 8591 8186
rect 8557 8099 8591 8101
rect 8557 8063 8591 8065
rect 8557 7978 8591 7997
rect 8671 8149 8705 8183
rect 8671 8081 8705 8115
rect 8671 8013 8705 8047
rect 8671 7945 8705 7979
rect 6895 7833 6929 7911
rect 7055 7901 7102 7935
rect 7138 7901 7172 7935
rect 7208 7901 7255 7935
rect 8345 7901 8392 7935
rect 8428 7901 8462 7935
rect 8498 7901 8545 7935
rect 8671 7833 8705 7911
rect 6895 7799 7015 7833
rect 7049 7799 7083 7833
rect 7117 7799 7151 7833
rect 7185 7799 7219 7833
rect 7253 7799 7287 7833
rect 7321 7799 7355 7833
rect 7389 7799 7423 7833
rect 7457 7799 7491 7833
rect 7525 7799 7559 7833
rect 7593 7799 7627 7833
rect 7661 7799 7695 7833
rect 7729 7799 7763 7833
rect 7797 7799 7831 7833
rect 7865 7799 7899 7833
rect 7933 7799 7967 7833
rect 8001 7799 8035 7833
rect 8069 7799 8103 7833
rect 8137 7799 8171 7833
rect 8205 7799 8239 7833
rect 8273 7799 8307 7833
rect 8341 7799 8375 7833
rect 8409 7799 8443 7833
rect 8477 7799 8511 7833
rect 8545 7799 8579 7833
rect 8613 7799 8705 7833
rect 1518 7730 1552 7764
rect -2322 7662 -2288 7696
rect -2162 7678 -2115 7712
rect -2079 7678 -2045 7712
rect -2009 7678 -1962 7712
rect 1192 7678 1239 7712
rect 1275 7678 1309 7712
rect 1345 7678 1392 7712
rect -2322 7594 -2288 7628
rect 1518 7662 1552 7696
rect -2162 7570 -2115 7604
rect -2079 7570 -2045 7604
rect -2009 7570 -1962 7604
rect -1904 7570 -1857 7604
rect -1821 7570 -1787 7604
rect -1751 7570 -1704 7604
rect -1646 7570 -1599 7604
rect -1563 7570 -1529 7604
rect -1493 7570 -1446 7604
rect -1388 7570 -1341 7604
rect -1305 7570 -1271 7604
rect -1235 7570 -1188 7604
rect -1130 7570 -1083 7604
rect -1047 7570 -1013 7604
rect -977 7570 -930 7604
rect -356 7570 -309 7604
rect -273 7570 -239 7604
rect -203 7570 -156 7604
rect -98 7570 -51 7604
rect -15 7570 19 7604
rect 55 7570 102 7604
rect 676 7570 723 7604
rect 759 7570 793 7604
rect 829 7570 876 7604
rect 934 7570 981 7604
rect 1017 7570 1051 7604
rect 1087 7570 1134 7604
rect 1192 7570 1239 7604
rect 1275 7570 1309 7604
rect 1345 7570 1392 7604
rect 1518 7594 1552 7628
rect -2322 7526 -2288 7560
rect -2322 7458 -2288 7492
rect -2322 7390 -2288 7424
rect -2322 7322 -2288 7356
rect -2208 7517 -2174 7536
rect -2208 7449 -2174 7451
rect -2208 7413 -2174 7415
rect -2208 7328 -2174 7347
rect -1950 7517 -1916 7536
rect -1950 7449 -1916 7451
rect -1950 7413 -1916 7415
rect -1950 7328 -1916 7347
rect -1692 7517 -1658 7536
rect -1692 7449 -1658 7451
rect -1692 7413 -1658 7415
rect -1692 7328 -1658 7347
rect -1434 7517 -1400 7536
rect -1434 7449 -1400 7451
rect -1434 7413 -1400 7415
rect -1434 7328 -1400 7347
rect -1176 7517 -1142 7536
rect -1176 7449 -1142 7451
rect -1176 7413 -1142 7415
rect -1176 7328 -1142 7347
rect -918 7517 -884 7536
rect -918 7449 -884 7451
rect -918 7413 -884 7415
rect -918 7328 -884 7347
rect -660 7517 -626 7536
rect -660 7449 -626 7451
rect -660 7413 -626 7415
rect -660 7328 -626 7347
rect -402 7517 -368 7536
rect -402 7449 -368 7451
rect -402 7413 -368 7415
rect -402 7328 -368 7347
rect -144 7517 -110 7536
rect -144 7449 -110 7451
rect -144 7413 -110 7415
rect -144 7328 -110 7347
rect 114 7517 148 7536
rect 114 7449 148 7451
rect 114 7413 148 7415
rect 114 7328 148 7347
rect 372 7517 406 7536
rect 372 7449 406 7451
rect 372 7413 406 7415
rect 372 7328 406 7347
rect 630 7517 664 7536
rect 630 7449 664 7451
rect 630 7413 664 7415
rect 630 7328 664 7347
rect 888 7517 922 7536
rect 888 7449 922 7451
rect 888 7413 922 7415
rect 888 7328 922 7347
rect 1146 7517 1180 7536
rect 1146 7449 1180 7451
rect 1146 7413 1180 7415
rect 1146 7328 1180 7347
rect 1404 7517 1438 7536
rect 1404 7449 1438 7451
rect 1404 7413 1438 7415
rect 1404 7328 1438 7347
rect 1518 7526 1552 7560
rect 1518 7458 1552 7492
rect 9741 7605 10350 7761
rect 9741 7603 9940 7605
rect 10262 7603 10350 7605
rect 9741 7501 9914 7603
rect 10288 7501 10350 7603
rect 9741 7499 9940 7501
rect 10262 7499 10350 7501
rect 1518 7390 1552 7424
rect 1518 7322 1552 7356
rect -2322 7254 -2288 7288
rect -2162 7260 -2115 7294
rect -2079 7260 -2045 7294
rect -2009 7260 -1962 7294
rect -872 7260 -825 7294
rect -789 7260 -755 7294
rect -719 7260 -672 7294
rect -614 7260 -567 7294
rect -531 7260 -497 7294
rect -461 7260 -414 7294
rect 160 7260 207 7294
rect 243 7260 277 7294
rect 313 7260 360 7294
rect 418 7260 465 7294
rect 501 7260 535 7294
rect 571 7260 618 7294
rect 1192 7260 1239 7294
rect 1275 7260 1309 7294
rect 1345 7260 1392 7294
rect -2322 7186 -2288 7220
rect 1518 7254 1552 7288
rect 1518 7186 1552 7220
rect -2162 7152 -2115 7186
rect -2079 7152 -2045 7186
rect -2009 7152 -1962 7186
rect -1904 7152 -1857 7186
rect -1821 7152 -1787 7186
rect -1751 7152 -1704 7186
rect -1646 7152 -1599 7186
rect -1563 7152 -1529 7186
rect -1493 7152 -1446 7186
rect -872 7152 -825 7186
rect -789 7152 -755 7186
rect -719 7152 -672 7186
rect -614 7152 -567 7186
rect -531 7152 -497 7186
rect -461 7152 -414 7186
rect 160 7152 207 7186
rect 243 7152 277 7186
rect 313 7152 360 7186
rect 418 7152 465 7186
rect 501 7152 535 7186
rect 571 7152 618 7186
rect 1192 7152 1239 7186
rect 1275 7152 1309 7186
rect 1345 7152 1392 7186
rect -2322 7118 -2288 7152
rect 1518 7118 1552 7152
rect -2322 7050 -2288 7084
rect -2322 6982 -2288 7016
rect -2322 6914 -2288 6948
rect -2208 7099 -2174 7118
rect -2208 7031 -2174 7033
rect -2208 6995 -2174 6997
rect -2208 6910 -2174 6929
rect -1950 7099 -1916 7118
rect -1950 7031 -1916 7033
rect -1950 6995 -1916 6997
rect -1950 6910 -1916 6929
rect -1692 7099 -1658 7118
rect -1692 7031 -1658 7033
rect -1692 6995 -1658 6997
rect -1692 6910 -1658 6929
rect -1434 7099 -1400 7118
rect -1434 7031 -1400 7033
rect -1434 6995 -1400 6997
rect -1434 6910 -1400 6929
rect -1176 7099 -1142 7118
rect -1176 7031 -1142 7033
rect -1176 6995 -1142 6997
rect -1176 6910 -1142 6929
rect -918 7099 -884 7118
rect -918 7031 -884 7033
rect -918 6995 -884 6997
rect -918 6910 -884 6929
rect -660 7099 -626 7118
rect -660 7031 -626 7033
rect -660 6995 -626 6997
rect -660 6910 -626 6929
rect -402 7099 -368 7118
rect -402 7031 -368 7033
rect -402 6995 -368 6997
rect -402 6910 -368 6929
rect -144 7099 -110 7118
rect -144 7031 -110 7033
rect -144 6995 -110 6997
rect -144 6910 -110 6929
rect 114 7099 148 7118
rect 114 7031 148 7033
rect 114 6995 148 6997
rect 114 6910 148 6929
rect 372 7099 406 7118
rect 372 7031 406 7033
rect 372 6995 406 6997
rect 372 6910 406 6929
rect 630 7099 664 7118
rect 630 7031 664 7033
rect 630 6995 664 6997
rect 630 6910 664 6929
rect 888 7099 922 7118
rect 888 7031 922 7033
rect 888 6995 922 6997
rect 888 6910 922 6929
rect 1146 7099 1180 7118
rect 1146 7031 1180 7033
rect 1146 6995 1180 6997
rect 1146 6910 1180 6929
rect 1404 7099 1438 7118
rect 1404 7031 1438 7033
rect 1404 6995 1438 6997
rect 1404 6910 1438 6929
rect 1518 7050 1552 7084
rect 1518 6982 1552 7016
rect 1518 6914 1552 6948
rect -2322 6846 -2288 6880
rect -2162 6842 -2115 6876
rect -2079 6842 -2045 6876
rect -2009 6842 -1962 6876
rect -1388 6842 -1341 6876
rect -1305 6842 -1271 6876
rect -1235 6842 -1188 6876
rect -1130 6842 -1083 6876
rect -1047 6842 -1013 6876
rect -977 6842 -930 6876
rect -356 6842 -309 6876
rect -273 6842 -239 6876
rect -203 6842 -156 6876
rect -98 6842 -51 6876
rect -15 6842 19 6876
rect 55 6842 102 6876
rect 676 6842 723 6876
rect 759 6842 793 6876
rect 829 6842 876 6876
rect 934 6842 981 6876
rect 1017 6842 1051 6876
rect 1087 6842 1134 6876
rect 1192 6842 1239 6876
rect 1275 6842 1309 6876
rect 1345 6842 1392 6876
rect 1518 6846 1552 6880
rect -2322 6778 -2288 6812
rect 1518 6778 1552 6812
rect -2322 6710 -2288 6744
rect -2162 6734 -2115 6768
rect -2079 6734 -2045 6768
rect -2009 6734 -1962 6768
rect -1388 6734 -1341 6768
rect -1305 6734 -1271 6768
rect -1235 6734 -1188 6768
rect -1130 6734 -1083 6768
rect -1047 6734 -1013 6768
rect -977 6734 -930 6768
rect -356 6734 -309 6768
rect -273 6734 -239 6768
rect -203 6734 -156 6768
rect -98 6734 -51 6768
rect -15 6734 19 6768
rect 55 6734 102 6768
rect 676 6734 723 6768
rect 759 6734 793 6768
rect 829 6734 876 6768
rect 934 6734 981 6768
rect 1017 6734 1051 6768
rect 1087 6734 1134 6768
rect 1192 6734 1239 6768
rect 1275 6734 1309 6768
rect 1345 6734 1392 6768
rect 1518 6710 1552 6744
rect -2322 6642 -2288 6676
rect -2322 6574 -2288 6608
rect -2322 6506 -2288 6540
rect -2208 6681 -2174 6700
rect -2208 6613 -2174 6615
rect -2208 6577 -2174 6579
rect -2208 6492 -2174 6511
rect -1950 6681 -1916 6700
rect -1950 6613 -1916 6615
rect -1950 6577 -1916 6579
rect -1950 6492 -1916 6511
rect -1692 6681 -1658 6700
rect -1692 6613 -1658 6615
rect -1692 6577 -1658 6579
rect -1692 6492 -1658 6511
rect -1434 6681 -1400 6700
rect -1434 6613 -1400 6615
rect -1434 6577 -1400 6579
rect -1434 6492 -1400 6511
rect -1176 6681 -1142 6700
rect -1176 6613 -1142 6615
rect -1176 6577 -1142 6579
rect -1176 6492 -1142 6511
rect -918 6681 -884 6700
rect -918 6613 -884 6615
rect -918 6577 -884 6579
rect -918 6492 -884 6511
rect -660 6681 -626 6700
rect -660 6613 -626 6615
rect -660 6577 -626 6579
rect -660 6492 -626 6511
rect -402 6681 -368 6700
rect -402 6613 -368 6615
rect -402 6577 -368 6579
rect -402 6492 -368 6511
rect -144 6681 -110 6700
rect -144 6613 -110 6615
rect -144 6577 -110 6579
rect -144 6492 -110 6511
rect 114 6681 148 6700
rect 114 6613 148 6615
rect 114 6577 148 6579
rect 114 6492 148 6511
rect 372 6681 406 6700
rect 372 6613 406 6615
rect 372 6577 406 6579
rect 372 6492 406 6511
rect 630 6681 664 6700
rect 630 6613 664 6615
rect 630 6577 664 6579
rect 630 6492 664 6511
rect 888 6681 922 6700
rect 888 6613 922 6615
rect 888 6577 922 6579
rect 888 6492 922 6511
rect 1146 6681 1180 6700
rect 1146 6613 1180 6615
rect 1146 6577 1180 6579
rect 1146 6492 1180 6511
rect 1404 6681 1438 6700
rect 1404 6613 1438 6615
rect 1404 6577 1438 6579
rect 1404 6492 1438 6511
rect 1518 6642 1552 6676
rect 1518 6574 1552 6608
rect 1518 6506 1552 6540
rect -2322 6438 -2288 6472
rect -2162 6424 -2115 6458
rect -2079 6424 -2045 6458
rect -2009 6424 -1962 6458
rect -1904 6424 -1857 6458
rect -1821 6424 -1787 6458
rect -1751 6424 -1704 6458
rect -1646 6424 -1599 6458
rect -1563 6424 -1529 6458
rect -1493 6424 -1446 6458
rect -872 6424 -825 6458
rect -789 6424 -755 6458
rect -719 6424 -672 6458
rect -614 6424 -567 6458
rect -531 6424 -497 6458
rect -461 6424 -414 6458
rect 160 6424 207 6458
rect 243 6424 277 6458
rect 313 6424 360 6458
rect 418 6424 465 6458
rect 501 6424 535 6458
rect 571 6424 618 6458
rect 1192 6424 1239 6458
rect 1275 6424 1309 6458
rect 1345 6424 1392 6458
rect 1518 6438 1552 6472
rect -2322 6370 -2288 6404
rect 1518 6370 1552 6404
rect -2322 6302 -2288 6336
rect -2162 6316 -2115 6350
rect -2079 6316 -2045 6350
rect -2009 6316 -1962 6350
rect -1904 6316 -1857 6350
rect -1821 6316 -1787 6350
rect -1751 6316 -1704 6350
rect -1646 6316 -1599 6350
rect -1563 6316 -1529 6350
rect -1493 6316 -1446 6350
rect -872 6316 -825 6350
rect -789 6316 -755 6350
rect -719 6316 -672 6350
rect -614 6316 -567 6350
rect -531 6316 -497 6350
rect -461 6316 -414 6350
rect 160 6316 207 6350
rect 243 6316 277 6350
rect 313 6316 360 6350
rect 418 6316 465 6350
rect 501 6316 535 6350
rect 571 6316 618 6350
rect 1192 6316 1239 6350
rect 1275 6316 1309 6350
rect 1345 6316 1392 6350
rect 1518 6302 1552 6336
rect -2322 6234 -2288 6268
rect -2322 6166 -2288 6200
rect -2322 6098 -2288 6132
rect -2208 6263 -2174 6282
rect -2208 6195 -2174 6197
rect -2208 6159 -2174 6161
rect -2208 6074 -2174 6093
rect -1950 6263 -1916 6282
rect -1950 6195 -1916 6197
rect -1950 6159 -1916 6161
rect -1950 6074 -1916 6093
rect -1692 6263 -1658 6282
rect -1692 6195 -1658 6197
rect -1692 6159 -1658 6161
rect -1692 6074 -1658 6093
rect -1434 6263 -1400 6282
rect -1434 6195 -1400 6197
rect -1434 6159 -1400 6161
rect -1434 6074 -1400 6093
rect -1176 6263 -1142 6282
rect -1176 6195 -1142 6197
rect -1176 6159 -1142 6161
rect -1176 6074 -1142 6093
rect -918 6263 -884 6282
rect -918 6195 -884 6197
rect -918 6159 -884 6161
rect -918 6074 -884 6093
rect -660 6263 -626 6282
rect -660 6195 -626 6197
rect -660 6159 -626 6161
rect -660 6074 -626 6093
rect -402 6263 -368 6282
rect -402 6195 -368 6197
rect -402 6159 -368 6161
rect -402 6074 -368 6093
rect -144 6263 -110 6282
rect -144 6195 -110 6197
rect -144 6159 -110 6161
rect -144 6074 -110 6093
rect 114 6263 148 6282
rect 114 6195 148 6197
rect 114 6159 148 6161
rect 114 6074 148 6093
rect 372 6263 406 6282
rect 372 6195 406 6197
rect 372 6159 406 6161
rect 372 6074 406 6093
rect 630 6263 664 6282
rect 630 6195 664 6197
rect 630 6159 664 6161
rect 630 6074 664 6093
rect 888 6263 922 6282
rect 888 6195 922 6197
rect 888 6159 922 6161
rect 888 6074 922 6093
rect 1146 6263 1180 6282
rect 1146 6195 1180 6197
rect 1146 6159 1180 6161
rect 1146 6074 1180 6093
rect 1404 6263 1438 6282
rect 1404 6195 1438 6197
rect 1404 6159 1438 6161
rect 1404 6074 1438 6093
rect 1518 6234 1552 6268
rect 1518 6166 1552 6200
rect 1518 6098 1552 6132
rect -2322 6030 -2288 6064
rect -2162 6006 -2115 6040
rect -2079 6006 -2045 6040
rect -2009 6006 -1962 6040
rect -1388 6006 -1341 6040
rect -1305 6006 -1271 6040
rect -1235 6006 -1188 6040
rect -1130 6006 -1083 6040
rect -1047 6006 -1013 6040
rect -977 6006 -930 6040
rect -356 6006 -309 6040
rect -273 6006 -239 6040
rect -203 6006 -156 6040
rect -98 6006 -51 6040
rect -15 6006 19 6040
rect 55 6006 102 6040
rect 676 6006 723 6040
rect 759 6006 793 6040
rect 829 6006 876 6040
rect 934 6006 981 6040
rect 1017 6006 1051 6040
rect 1087 6006 1134 6040
rect 1192 6006 1239 6040
rect 1275 6006 1309 6040
rect 1345 6006 1392 6040
rect 1518 6030 1552 6064
rect -2322 5962 -2288 5996
rect 1518 5962 1552 5996
rect -2322 5894 -2288 5928
rect -2162 5898 -2115 5932
rect -2079 5898 -2045 5932
rect -2009 5898 -1962 5932
rect -1388 5898 -1341 5932
rect -1305 5898 -1271 5932
rect -1235 5898 -1188 5932
rect -1130 5898 -1083 5932
rect -1047 5898 -1013 5932
rect -977 5898 -930 5932
rect -356 5898 -309 5932
rect -273 5898 -239 5932
rect -203 5898 -156 5932
rect -98 5898 -51 5932
rect -15 5898 19 5932
rect 55 5898 102 5932
rect 676 5898 723 5932
rect 759 5898 793 5932
rect 829 5898 876 5932
rect 934 5898 981 5932
rect 1017 5898 1051 5932
rect 1087 5898 1134 5932
rect 1192 5898 1239 5932
rect 1275 5898 1309 5932
rect 1345 5898 1392 5932
rect 1518 5894 1552 5928
rect -2322 5826 -2288 5860
rect -2322 5758 -2288 5792
rect -2322 5690 -2288 5724
rect -2208 5845 -2174 5864
rect -2208 5777 -2174 5779
rect -2208 5741 -2174 5743
rect -2208 5656 -2174 5675
rect -1950 5845 -1916 5864
rect -1950 5777 -1916 5779
rect -1950 5741 -1916 5743
rect -1950 5656 -1916 5675
rect -1692 5845 -1658 5864
rect -1692 5777 -1658 5779
rect -1692 5741 -1658 5743
rect -1692 5656 -1658 5675
rect -1434 5845 -1400 5864
rect -1434 5777 -1400 5779
rect -1434 5741 -1400 5743
rect -1434 5656 -1400 5675
rect -1176 5845 -1142 5864
rect -1176 5777 -1142 5779
rect -1176 5741 -1142 5743
rect -1176 5656 -1142 5675
rect -918 5845 -884 5864
rect -918 5777 -884 5779
rect -918 5741 -884 5743
rect -918 5656 -884 5675
rect -660 5845 -626 5864
rect -660 5777 -626 5779
rect -660 5741 -626 5743
rect -660 5656 -626 5675
rect -402 5845 -368 5864
rect -402 5777 -368 5779
rect -402 5741 -368 5743
rect -402 5656 -368 5675
rect -144 5845 -110 5864
rect -144 5777 -110 5779
rect -144 5741 -110 5743
rect -144 5656 -110 5675
rect 114 5845 148 5864
rect 114 5777 148 5779
rect 114 5741 148 5743
rect 114 5656 148 5675
rect 372 5845 406 5864
rect 372 5777 406 5779
rect 372 5741 406 5743
rect 372 5656 406 5675
rect 630 5845 664 5864
rect 630 5777 664 5779
rect 630 5741 664 5743
rect 630 5656 664 5675
rect 888 5845 922 5864
rect 888 5777 922 5779
rect 888 5741 922 5743
rect 888 5656 922 5675
rect 1146 5845 1180 5864
rect 1146 5777 1180 5779
rect 1146 5741 1180 5743
rect 1146 5656 1180 5675
rect 1404 5845 1438 5864
rect 1404 5777 1438 5779
rect 1404 5741 1438 5743
rect 1404 5656 1438 5675
rect 1518 5826 1552 5860
rect 1518 5758 1552 5792
rect 1518 5690 1552 5724
rect -2322 5622 -2288 5656
rect 1518 5622 1552 5656
rect -2162 5588 -2115 5622
rect -2079 5588 -2045 5622
rect -2009 5588 -1962 5622
rect -1904 5588 -1857 5622
rect -1821 5588 -1787 5622
rect -1751 5588 -1704 5622
rect -1646 5588 -1599 5622
rect -1563 5588 -1529 5622
rect -1493 5588 -1446 5622
rect -872 5588 -825 5622
rect -789 5588 -755 5622
rect -719 5588 -672 5622
rect -614 5588 -567 5622
rect -531 5588 -497 5622
rect -461 5588 -414 5622
rect 160 5588 207 5622
rect 243 5588 277 5622
rect 313 5588 360 5622
rect 418 5588 465 5622
rect 501 5588 535 5622
rect 571 5588 618 5622
rect 1192 5588 1239 5622
rect 1275 5588 1309 5622
rect 1345 5588 1392 5622
rect -2322 5554 -2288 5588
rect -2322 5486 -2288 5520
rect 1518 5554 1552 5588
rect -2162 5480 -2115 5514
rect -2079 5480 -2045 5514
rect -2009 5480 -1962 5514
rect -1904 5480 -1857 5514
rect -1821 5480 -1787 5514
rect -1751 5480 -1704 5514
rect -1646 5480 -1599 5514
rect -1563 5480 -1529 5514
rect -1493 5480 -1446 5514
rect -872 5480 -825 5514
rect -789 5480 -755 5514
rect -719 5480 -672 5514
rect -614 5480 -567 5514
rect -531 5480 -497 5514
rect -461 5480 -414 5514
rect 160 5480 207 5514
rect 243 5480 277 5514
rect 313 5480 360 5514
rect 418 5480 465 5514
rect 501 5480 535 5514
rect 571 5480 618 5514
rect 1192 5480 1239 5514
rect 1275 5480 1309 5514
rect 1345 5480 1392 5514
rect 1518 5486 1552 5520
rect -2322 5418 -2288 5452
rect -2322 5350 -2288 5384
rect -2322 5282 -2288 5316
rect -2322 5214 -2288 5248
rect -2208 5427 -2174 5446
rect -2208 5359 -2174 5361
rect -2208 5323 -2174 5325
rect -2208 5238 -2174 5257
rect -1950 5427 -1916 5446
rect -1950 5359 -1916 5361
rect -1950 5323 -1916 5325
rect -1950 5238 -1916 5257
rect -1692 5427 -1658 5446
rect -1692 5359 -1658 5361
rect -1692 5323 -1658 5325
rect -1692 5238 -1658 5257
rect -1434 5427 -1400 5446
rect -1434 5359 -1400 5361
rect -1434 5323 -1400 5325
rect -1434 5238 -1400 5257
rect -1176 5427 -1142 5446
rect -1176 5359 -1142 5361
rect -1176 5323 -1142 5325
rect -1176 5238 -1142 5257
rect -918 5427 -884 5446
rect -918 5359 -884 5361
rect -918 5323 -884 5325
rect -918 5238 -884 5257
rect -660 5427 -626 5446
rect -660 5359 -626 5361
rect -660 5323 -626 5325
rect -660 5238 -626 5257
rect -402 5427 -368 5446
rect -402 5359 -368 5361
rect -402 5323 -368 5325
rect -402 5238 -368 5257
rect -144 5427 -110 5446
rect -144 5359 -110 5361
rect -144 5323 -110 5325
rect -144 5238 -110 5257
rect 114 5427 148 5446
rect 114 5359 148 5361
rect 114 5323 148 5325
rect 114 5238 148 5257
rect 372 5427 406 5446
rect 372 5359 406 5361
rect 372 5323 406 5325
rect 372 5238 406 5257
rect 630 5427 664 5446
rect 630 5359 664 5361
rect 630 5323 664 5325
rect 630 5238 664 5257
rect 888 5427 922 5446
rect 888 5359 922 5361
rect 888 5323 922 5325
rect 888 5238 922 5257
rect 1146 5427 1180 5446
rect 1146 5359 1180 5361
rect 1146 5323 1180 5325
rect 1146 5238 1180 5257
rect 1404 5427 1438 5446
rect 1404 5359 1438 5361
rect 1404 5323 1438 5325
rect 1404 5238 1438 5257
rect 1518 5418 1552 5452
rect 1518 5350 1552 5384
rect 1518 5282 1552 5316
rect 1518 5214 1552 5248
rect -2322 5146 -2288 5180
rect -2162 5170 -2115 5204
rect -2079 5170 -2045 5204
rect -2009 5170 -1962 5204
rect -1388 5170 -1341 5204
rect -1305 5170 -1271 5204
rect -1235 5170 -1188 5204
rect -1130 5170 -1083 5204
rect -1047 5170 -1013 5204
rect -977 5170 -930 5204
rect -356 5170 -309 5204
rect -273 5170 -239 5204
rect -203 5170 -156 5204
rect -98 5170 -51 5204
rect -15 5170 19 5204
rect 55 5170 102 5204
rect 676 5170 723 5204
rect 759 5170 793 5204
rect 829 5170 876 5204
rect 934 5170 981 5204
rect 1017 5170 1051 5204
rect 1087 5170 1134 5204
rect 1192 5170 1239 5204
rect 1275 5170 1309 5204
rect 1345 5170 1392 5204
rect -2322 5078 -2288 5112
rect 1518 5146 1552 5180
rect -2162 5062 -2115 5096
rect -2079 5062 -2045 5096
rect -2009 5062 -1962 5096
rect -1388 5062 -1341 5096
rect -1305 5062 -1271 5096
rect -1235 5062 -1188 5096
rect -1130 5062 -1083 5096
rect -1047 5062 -1013 5096
rect -977 5062 -930 5096
rect -356 5062 -309 5096
rect -273 5062 -239 5096
rect -203 5062 -156 5096
rect -98 5062 -51 5096
rect -15 5062 19 5096
rect 55 5062 102 5096
rect 676 5062 723 5096
rect 759 5062 793 5096
rect 829 5062 876 5096
rect 934 5062 981 5096
rect 1017 5062 1051 5096
rect 1087 5062 1134 5096
rect 1192 5062 1239 5096
rect 1275 5062 1309 5096
rect 1345 5062 1392 5096
rect 1518 5078 1552 5112
rect -2322 5010 -2288 5044
rect -2322 4942 -2288 4976
rect -2322 4874 -2288 4908
rect -2322 4806 -2288 4840
rect -2208 5009 -2174 5028
rect -2208 4941 -2174 4943
rect -2208 4905 -2174 4907
rect -2208 4820 -2174 4839
rect -1950 5009 -1916 5028
rect -1950 4941 -1916 4943
rect -1950 4905 -1916 4907
rect -1950 4820 -1916 4839
rect -1692 5009 -1658 5028
rect -1692 4941 -1658 4943
rect -1692 4905 -1658 4907
rect -1692 4820 -1658 4839
rect -1434 5009 -1400 5028
rect -1434 4941 -1400 4943
rect -1434 4905 -1400 4907
rect -1434 4820 -1400 4839
rect -1176 5009 -1142 5028
rect -1176 4941 -1142 4943
rect -1176 4905 -1142 4907
rect -1176 4820 -1142 4839
rect -918 5009 -884 5028
rect -918 4941 -884 4943
rect -918 4905 -884 4907
rect -918 4820 -884 4839
rect -660 5009 -626 5028
rect -660 4941 -626 4943
rect -660 4905 -626 4907
rect -660 4820 -626 4839
rect -402 5009 -368 5028
rect -402 4941 -368 4943
rect -402 4905 -368 4907
rect -402 4820 -368 4839
rect -144 5009 -110 5028
rect -144 4941 -110 4943
rect -144 4905 -110 4907
rect -144 4820 -110 4839
rect 114 5009 148 5028
rect 114 4941 148 4943
rect 114 4905 148 4907
rect 114 4820 148 4839
rect 372 5009 406 5028
rect 372 4941 406 4943
rect 372 4905 406 4907
rect 372 4820 406 4839
rect 630 5009 664 5028
rect 630 4941 664 4943
rect 630 4905 664 4907
rect 630 4820 664 4839
rect 888 5009 922 5028
rect 888 4941 922 4943
rect 888 4905 922 4907
rect 888 4820 922 4839
rect 1146 5009 1180 5028
rect 1146 4941 1180 4943
rect 1146 4905 1180 4907
rect 1146 4820 1180 4839
rect 1404 5009 1438 5028
rect 1404 4941 1438 4943
rect 1404 4905 1438 4907
rect 1404 4820 1438 4839
rect 1518 5010 1552 5044
rect 1518 4942 1552 4976
rect 1518 4874 1552 4908
rect 1518 4806 1552 4840
rect -2322 4738 -2288 4772
rect -2162 4752 -2115 4786
rect -2079 4752 -2045 4786
rect -2009 4752 -1962 4786
rect -1904 4752 -1857 4786
rect -1821 4752 -1787 4786
rect -1751 4752 -1704 4786
rect -1646 4752 -1599 4786
rect -1563 4752 -1529 4786
rect -1493 4752 -1446 4786
rect -872 4752 -825 4786
rect -789 4752 -755 4786
rect -719 4752 -672 4786
rect -614 4752 -567 4786
rect -531 4752 -497 4786
rect -461 4752 -414 4786
rect 160 4752 207 4786
rect 243 4752 277 4786
rect 313 4752 360 4786
rect 418 4752 465 4786
rect 501 4752 535 4786
rect 571 4752 618 4786
rect 1192 4752 1239 4786
rect 1275 4752 1309 4786
rect 1345 4752 1392 4786
rect -2322 4670 -2288 4704
rect 1518 4738 1552 4772
rect -2162 4644 -2115 4678
rect -2079 4644 -2045 4678
rect -2009 4644 -1962 4678
rect -1904 4644 -1857 4678
rect -1821 4644 -1787 4678
rect -1751 4644 -1704 4678
rect -1646 4644 -1599 4678
rect -1563 4644 -1529 4678
rect -1493 4644 -1446 4678
rect -872 4644 -825 4678
rect -789 4644 -755 4678
rect -719 4644 -672 4678
rect -614 4644 -567 4678
rect -531 4644 -497 4678
rect -461 4644 -414 4678
rect 160 4644 207 4678
rect 243 4644 277 4678
rect 313 4644 360 4678
rect 418 4644 465 4678
rect 501 4644 535 4678
rect 571 4644 618 4678
rect 676 4644 723 4678
rect 759 4644 793 4678
rect 829 4644 876 4678
rect 934 4644 981 4678
rect 1017 4644 1051 4678
rect 1087 4644 1134 4678
rect 1192 4644 1239 4678
rect 1275 4644 1309 4678
rect 1345 4644 1392 4678
rect 1518 4670 1552 4704
rect -2322 4602 -2288 4636
rect -2322 4534 -2288 4568
rect -2322 4466 -2288 4500
rect -2322 4398 -2288 4432
rect -2208 4591 -2174 4610
rect -2208 4523 -2174 4525
rect -2208 4487 -2174 4489
rect -2208 4402 -2174 4421
rect -1950 4591 -1916 4610
rect -1950 4523 -1916 4525
rect -1950 4487 -1916 4489
rect -1950 4402 -1916 4421
rect -1692 4591 -1658 4610
rect -1692 4523 -1658 4525
rect -1692 4487 -1658 4489
rect -1692 4402 -1658 4421
rect -1434 4591 -1400 4610
rect -1434 4523 -1400 4525
rect -1434 4487 -1400 4489
rect -1434 4402 -1400 4421
rect -1176 4591 -1142 4610
rect -1176 4523 -1142 4525
rect -1176 4487 -1142 4489
rect -1176 4402 -1142 4421
rect -918 4591 -884 4610
rect -918 4523 -884 4525
rect -918 4487 -884 4489
rect -918 4402 -884 4421
rect -660 4591 -626 4610
rect -660 4523 -626 4525
rect -660 4487 -626 4489
rect -660 4402 -626 4421
rect -402 4591 -368 4610
rect -402 4523 -368 4525
rect -402 4487 -368 4489
rect -402 4402 -368 4421
rect -144 4591 -110 4610
rect -144 4523 -110 4525
rect -144 4487 -110 4489
rect -144 4402 -110 4421
rect 114 4591 148 4610
rect 114 4523 148 4525
rect 114 4487 148 4489
rect 114 4402 148 4421
rect 372 4591 406 4610
rect 372 4523 406 4525
rect 372 4487 406 4489
rect 372 4402 406 4421
rect 630 4591 664 4610
rect 630 4523 664 4525
rect 630 4487 664 4489
rect 630 4402 664 4421
rect 888 4591 922 4610
rect 888 4523 922 4525
rect 888 4487 922 4489
rect 888 4402 922 4421
rect 1146 4591 1180 4610
rect 1146 4523 1180 4525
rect 1146 4487 1180 4489
rect 1146 4402 1180 4421
rect 1404 4591 1438 4610
rect 1404 4523 1438 4525
rect 1404 4487 1438 4489
rect 1404 4402 1438 4421
rect 1518 4602 1552 4636
rect 1518 4534 1552 4568
rect 1518 4466 1552 4500
rect 1518 4398 1552 4432
rect -2322 4330 -2288 4364
rect -2162 4334 -2115 4368
rect -2079 4334 -2045 4368
rect -2009 4334 -1962 4368
rect -1388 4334 -1341 4368
rect -1305 4334 -1271 4368
rect -1235 4334 -1188 4368
rect -1130 4334 -1083 4368
rect -1047 4334 -1013 4368
rect -977 4334 -930 4368
rect -356 4334 -309 4368
rect -273 4334 -239 4368
rect -203 4334 -156 4368
rect -98 4334 -51 4368
rect -15 4334 19 4368
rect 55 4334 102 4368
rect 1192 4334 1239 4368
rect 1275 4334 1309 4368
rect 1345 4334 1392 4368
rect -2322 4262 -2288 4296
rect 1518 4330 1552 4364
rect 1518 4262 1552 4296
rect -2322 4194 -2288 4228
rect -2162 4226 -2115 4260
rect -2079 4226 -2045 4260
rect -2009 4226 -1962 4260
rect -1904 4226 -1857 4260
rect -1821 4226 -1787 4260
rect -1751 4226 -1704 4260
rect -1646 4226 -1599 4260
rect -1563 4226 -1529 4260
rect -1493 4226 -1446 4260
rect -1388 4226 -1341 4260
rect -1305 4226 -1271 4260
rect -1235 4226 -1188 4260
rect -1130 4226 -1083 4260
rect -1047 4226 -1013 4260
rect -977 4226 -930 4260
rect -872 4226 -825 4260
rect -789 4226 -755 4260
rect -719 4226 -672 4260
rect -614 4226 -567 4260
rect -531 4226 -497 4260
rect -461 4226 -414 4260
rect -356 4226 -309 4260
rect -273 4226 -239 4260
rect -203 4226 -156 4260
rect -98 4226 -51 4260
rect -15 4226 19 4260
rect 55 4226 102 4260
rect 160 4226 207 4260
rect 243 4226 277 4260
rect 313 4226 360 4260
rect 418 4226 465 4260
rect 501 4226 535 4260
rect 571 4226 618 4260
rect 676 4226 723 4260
rect 759 4226 793 4260
rect 829 4226 876 4260
rect 934 4226 981 4260
rect 1017 4226 1051 4260
rect 1087 4226 1134 4260
rect 1192 4226 1239 4260
rect 1275 4226 1309 4260
rect 1345 4226 1392 4260
rect 1518 4194 1552 4228
rect -2322 4126 -2288 4160
rect -2322 4058 -2288 4092
rect -2322 3990 -2288 4024
rect -2208 4173 -2174 4192
rect -2208 4105 -2174 4107
rect -2208 4069 -2174 4071
rect -2208 3984 -2174 4003
rect -1950 4173 -1916 4192
rect -1950 4105 -1916 4107
rect -1950 4069 -1916 4071
rect -1950 3984 -1916 4003
rect -1692 4173 -1658 4192
rect -1692 4105 -1658 4107
rect -1692 4069 -1658 4071
rect -1692 3984 -1658 4003
rect -1434 4173 -1400 4192
rect -1434 4105 -1400 4107
rect -1434 4069 -1400 4071
rect -1434 3984 -1400 4003
rect -1176 4173 -1142 4192
rect -1176 4105 -1142 4107
rect -1176 4069 -1142 4071
rect -1176 3984 -1142 4003
rect -918 4173 -884 4192
rect -918 4105 -884 4107
rect -918 4069 -884 4071
rect -918 3984 -884 4003
rect -660 4173 -626 4192
rect -660 4105 -626 4107
rect -660 4069 -626 4071
rect -660 3984 -626 4003
rect -402 4173 -368 4192
rect -402 4105 -368 4107
rect -402 4069 -368 4071
rect -402 3984 -368 4003
rect -144 4173 -110 4192
rect -144 4105 -110 4107
rect -144 4069 -110 4071
rect -144 3984 -110 4003
rect 114 4173 148 4192
rect 114 4105 148 4107
rect 114 4069 148 4071
rect 114 3984 148 4003
rect 372 4173 406 4192
rect 372 4105 406 4107
rect 372 4069 406 4071
rect 372 3984 406 4003
rect 630 4173 664 4192
rect 630 4105 664 4107
rect 630 4069 664 4071
rect 630 3984 664 4003
rect 888 4173 922 4192
rect 888 4105 922 4107
rect 888 4069 922 4071
rect 888 3984 922 4003
rect 1146 4173 1180 4192
rect 1146 4105 1180 4107
rect 1146 4069 1180 4071
rect 1146 3984 1180 4003
rect 1404 4173 1438 4192
rect 1404 4105 1438 4107
rect 1404 4069 1438 4071
rect 1404 3984 1438 4003
rect 1518 4126 1552 4160
rect 1518 4058 1552 4092
rect 3508 7451 3628 7485
rect 3662 7451 3696 7485
rect 3730 7451 3764 7485
rect 3798 7451 3832 7485
rect 3866 7451 3900 7485
rect 3934 7451 3968 7485
rect 4002 7451 4036 7485
rect 4070 7451 4104 7485
rect 4138 7451 4172 7485
rect 4206 7451 4240 7485
rect 4274 7451 4308 7485
rect 4342 7451 4376 7485
rect 4410 7451 4444 7485
rect 4478 7451 4512 7485
rect 4546 7451 4580 7485
rect 4614 7451 4648 7485
rect 4682 7451 4716 7485
rect 4750 7451 4784 7485
rect 4818 7451 4852 7485
rect 4886 7451 4920 7485
rect 4954 7451 4988 7485
rect 5022 7451 5056 7485
rect 5090 7451 5124 7485
rect 5158 7451 5192 7485
rect 5226 7451 5260 7485
rect 5294 7451 5328 7485
rect 5362 7451 5396 7485
rect 5430 7451 5464 7485
rect 5498 7451 5532 7485
rect 5566 7451 5600 7485
rect 5634 7451 5668 7485
rect 5702 7451 5736 7485
rect 5770 7451 5804 7485
rect 5838 7451 5872 7485
rect 5906 7451 5940 7485
rect 5974 7451 6008 7485
rect 6042 7451 6076 7485
rect 6110 7451 6144 7485
rect 6178 7451 6212 7485
rect 6246 7451 6350 7485
rect 3508 7363 3542 7451
rect 3668 7349 3715 7383
rect 3751 7349 3785 7383
rect 3821 7349 3868 7383
rect 3926 7349 3973 7383
rect 4009 7349 4043 7383
rect 4079 7349 4126 7383
rect 4184 7349 4231 7383
rect 4267 7349 4301 7383
rect 4337 7349 4384 7383
rect 4442 7349 4489 7383
rect 4525 7349 4559 7383
rect 4595 7349 4642 7383
rect 4700 7349 4747 7383
rect 4783 7349 4817 7383
rect 4853 7349 4900 7383
rect 4958 7349 5005 7383
rect 5041 7349 5075 7383
rect 5111 7349 5158 7383
rect 5216 7349 5263 7383
rect 5299 7349 5333 7383
rect 5369 7349 5416 7383
rect 5474 7349 5521 7383
rect 5557 7349 5591 7383
rect 5627 7349 5674 7383
rect 5732 7349 5779 7383
rect 5815 7349 5849 7383
rect 5885 7349 5932 7383
rect 5990 7349 6037 7383
rect 6073 7349 6107 7383
rect 6143 7349 6190 7383
rect 6316 7363 6350 7451
rect 9741 7364 10350 7499
rect 3508 7295 3542 7329
rect 3508 7227 3542 7261
rect 3508 7159 3542 7193
rect 3508 7091 3542 7125
rect 3622 7296 3656 7315
rect 3622 7228 3656 7230
rect 3622 7192 3656 7194
rect 3622 7107 3656 7126
rect 3880 7296 3914 7315
rect 3880 7228 3914 7230
rect 3880 7192 3914 7194
rect 3880 7107 3914 7126
rect 4138 7296 4172 7315
rect 4138 7228 4172 7230
rect 4138 7192 4172 7194
rect 4138 7107 4172 7126
rect 4396 7296 4430 7315
rect 4396 7228 4430 7230
rect 4396 7192 4430 7194
rect 4396 7107 4430 7126
rect 4654 7296 4688 7315
rect 4654 7228 4688 7230
rect 4654 7192 4688 7194
rect 4654 7107 4688 7126
rect 4912 7296 4946 7315
rect 4912 7228 4946 7230
rect 4912 7192 4946 7194
rect 4912 7107 4946 7126
rect 5170 7296 5204 7315
rect 5170 7228 5204 7230
rect 5170 7192 5204 7194
rect 5170 7107 5204 7126
rect 5428 7296 5462 7315
rect 5428 7228 5462 7230
rect 5428 7192 5462 7194
rect 5428 7107 5462 7126
rect 5686 7296 5720 7315
rect 5686 7228 5720 7230
rect 5686 7192 5720 7194
rect 5686 7107 5720 7126
rect 5944 7296 5978 7315
rect 5944 7228 5978 7230
rect 5944 7192 5978 7194
rect 5944 7107 5978 7126
rect 6202 7296 6236 7315
rect 6202 7228 6236 7230
rect 6202 7192 6236 7194
rect 6202 7107 6236 7126
rect 6316 7295 6350 7329
rect 6316 7227 6350 7261
rect 6316 7159 6350 7193
rect 6316 7091 6350 7125
rect 3508 7023 3542 7057
rect 3668 7039 3715 7073
rect 3751 7039 3785 7073
rect 3821 7039 3868 7073
rect 5990 7039 6037 7073
rect 6073 7039 6107 7073
rect 6143 7039 6190 7073
rect 3508 6955 3542 6989
rect 6316 7023 6350 7057
rect 3668 6931 3715 6965
rect 3751 6931 3785 6965
rect 3821 6931 3868 6965
rect 3926 6931 3973 6965
rect 4009 6931 4043 6965
rect 4079 6931 4126 6965
rect 4184 6931 4231 6965
rect 4267 6931 4301 6965
rect 4337 6931 4384 6965
rect 4958 6931 5005 6965
rect 5041 6931 5075 6965
rect 5111 6931 5158 6965
rect 5216 6931 5263 6965
rect 5299 6931 5333 6965
rect 5369 6931 5416 6965
rect 5990 6931 6037 6965
rect 6073 6931 6107 6965
rect 6143 6931 6190 6965
rect 6316 6955 6350 6989
rect 3508 6887 3542 6921
rect 3508 6819 3542 6853
rect 3508 6751 3542 6785
rect 3508 6683 3542 6717
rect 3622 6878 3656 6897
rect 3622 6810 3656 6812
rect 3622 6774 3656 6776
rect 3622 6689 3656 6708
rect 3880 6878 3914 6897
rect 3880 6810 3914 6812
rect 3880 6774 3914 6776
rect 3880 6689 3914 6708
rect 4138 6878 4172 6897
rect 4138 6810 4172 6812
rect 4138 6774 4172 6776
rect 4138 6689 4172 6708
rect 4396 6878 4430 6897
rect 4396 6810 4430 6812
rect 4396 6774 4430 6776
rect 4396 6689 4430 6708
rect 4654 6878 4688 6897
rect 4654 6810 4688 6812
rect 4654 6774 4688 6776
rect 4654 6689 4688 6708
rect 4912 6878 4946 6897
rect 4912 6810 4946 6812
rect 4912 6774 4946 6776
rect 4912 6689 4946 6708
rect 5170 6878 5204 6897
rect 5170 6810 5204 6812
rect 5170 6774 5204 6776
rect 5170 6689 5204 6708
rect 5428 6878 5462 6897
rect 5428 6810 5462 6812
rect 5428 6774 5462 6776
rect 5428 6689 5462 6708
rect 5686 6878 5720 6897
rect 5686 6810 5720 6812
rect 5686 6774 5720 6776
rect 5686 6689 5720 6708
rect 5944 6878 5978 6897
rect 5944 6810 5978 6812
rect 5944 6774 5978 6776
rect 5944 6689 5978 6708
rect 6202 6878 6236 6897
rect 6202 6810 6236 6812
rect 6202 6774 6236 6776
rect 6202 6689 6236 6708
rect 6316 6887 6350 6921
rect 6316 6819 6350 6853
rect 6316 6751 6350 6785
rect 6316 6683 6350 6717
rect 3508 6615 3542 6649
rect 3668 6621 3715 6655
rect 3751 6621 3785 6655
rect 3821 6621 3868 6655
rect 4442 6621 4489 6655
rect 4525 6621 4559 6655
rect 4595 6621 4642 6655
rect 4700 6621 4747 6655
rect 4783 6621 4817 6655
rect 4853 6621 4900 6655
rect 5474 6621 5521 6655
rect 5557 6621 5591 6655
rect 5627 6621 5674 6655
rect 5732 6621 5779 6655
rect 5815 6621 5849 6655
rect 5885 6621 5932 6655
rect 5990 6621 6037 6655
rect 6073 6621 6107 6655
rect 6143 6621 6190 6655
rect 3508 6547 3542 6581
rect 6316 6615 6350 6649
rect 3668 6513 3715 6547
rect 3751 6513 3785 6547
rect 3821 6513 3868 6547
rect 4442 6513 4489 6547
rect 4525 6513 4559 6547
rect 4595 6513 4642 6547
rect 4700 6513 4747 6547
rect 4783 6513 4817 6547
rect 4853 6513 4900 6547
rect 5474 6513 5521 6547
rect 5557 6513 5591 6547
rect 5627 6513 5674 6547
rect 5732 6513 5779 6547
rect 5815 6513 5849 6547
rect 5885 6513 5932 6547
rect 5990 6513 6037 6547
rect 6073 6513 6107 6547
rect 6143 6513 6190 6547
rect 3508 6479 3542 6513
rect 6316 6479 6350 6581
rect 3508 6411 3542 6445
rect 3508 6343 3542 6377
rect 3508 6275 3542 6309
rect 3622 6460 3656 6479
rect 3622 6392 3656 6394
rect 3622 6356 3656 6358
rect 3622 6271 3656 6290
rect 3880 6460 3914 6479
rect 3880 6392 3914 6394
rect 3880 6356 3914 6358
rect 3880 6271 3914 6290
rect 4138 6460 4172 6479
rect 4138 6392 4172 6394
rect 4138 6356 4172 6358
rect 4138 6271 4172 6290
rect 4396 6460 4430 6479
rect 4396 6392 4430 6394
rect 4396 6356 4430 6358
rect 4396 6271 4430 6290
rect 4654 6460 4688 6479
rect 4654 6392 4688 6394
rect 4654 6356 4688 6358
rect 4654 6271 4688 6290
rect 4912 6460 4946 6479
rect 4912 6392 4946 6394
rect 4912 6356 4946 6358
rect 4912 6271 4946 6290
rect 5170 6460 5204 6479
rect 5170 6392 5204 6394
rect 5170 6356 5204 6358
rect 5170 6271 5204 6290
rect 5428 6460 5462 6479
rect 5428 6392 5462 6394
rect 5428 6356 5462 6358
rect 5428 6271 5462 6290
rect 5686 6460 5720 6479
rect 5686 6392 5720 6394
rect 5686 6356 5720 6358
rect 5686 6271 5720 6290
rect 5944 6460 5978 6479
rect 5944 6392 5978 6394
rect 5944 6356 5978 6358
rect 5944 6271 5978 6290
rect 6202 6460 6236 6479
rect 6202 6392 6236 6394
rect 6202 6356 6236 6358
rect 6202 6271 6236 6290
rect 6316 6411 6350 6445
rect 6316 6343 6350 6377
rect 6316 6275 6350 6309
rect 3508 6207 3542 6241
rect 3668 6203 3715 6237
rect 3751 6203 3785 6237
rect 3821 6203 3868 6237
rect 3926 6203 3973 6237
rect 4009 6203 4043 6237
rect 4079 6203 4126 6237
rect 4184 6203 4231 6237
rect 4267 6203 4301 6237
rect 4337 6203 4384 6237
rect 4958 6203 5005 6237
rect 5041 6203 5075 6237
rect 5111 6203 5158 6237
rect 5216 6203 5263 6237
rect 5299 6203 5333 6237
rect 5369 6203 5416 6237
rect 5990 6203 6037 6237
rect 6073 6203 6107 6237
rect 6143 6203 6190 6237
rect 6316 6207 6350 6241
rect 3508 6139 3542 6173
rect 6316 6139 6350 6173
rect 3508 6071 3542 6105
rect 3668 6095 3715 6129
rect 3751 6095 3785 6129
rect 3821 6095 3868 6129
rect 3926 6095 3973 6129
rect 4009 6095 4043 6129
rect 4079 6095 4126 6129
rect 4184 6095 4231 6129
rect 4267 6095 4301 6129
rect 4337 6095 4384 6129
rect 4958 6095 5005 6129
rect 5041 6095 5075 6129
rect 5111 6095 5158 6129
rect 5216 6095 5263 6129
rect 5299 6095 5333 6129
rect 5369 6095 5416 6129
rect 5990 6095 6037 6129
rect 6073 6095 6107 6129
rect 6143 6095 6190 6129
rect 6316 6071 6350 6105
rect 3508 6003 3542 6037
rect 3508 5935 3542 5969
rect 3508 5867 3542 5901
rect 3622 6042 3656 6061
rect 3622 5974 3656 5976
rect 3622 5938 3656 5940
rect 3622 5853 3656 5872
rect 3880 6042 3914 6061
rect 3880 5974 3914 5976
rect 3880 5938 3914 5940
rect 3880 5853 3914 5872
rect 4138 6042 4172 6061
rect 4138 5974 4172 5976
rect 4138 5938 4172 5940
rect 4138 5853 4172 5872
rect 4396 6042 4430 6061
rect 4396 5974 4430 5976
rect 4396 5938 4430 5940
rect 4396 5853 4430 5872
rect 4654 6042 4688 6061
rect 4654 5974 4688 5976
rect 4654 5938 4688 5940
rect 4654 5853 4688 5872
rect 4912 6042 4946 6061
rect 4912 5974 4946 5976
rect 4912 5938 4946 5940
rect 4912 5853 4946 5872
rect 5170 6042 5204 6061
rect 5170 5974 5204 5976
rect 5170 5938 5204 5940
rect 5170 5853 5204 5872
rect 5428 6042 5462 6061
rect 5428 5974 5462 5976
rect 5428 5938 5462 5940
rect 5428 5853 5462 5872
rect 5686 6042 5720 6061
rect 5686 5974 5720 5976
rect 5686 5938 5720 5940
rect 5686 5853 5720 5872
rect 5944 6042 5978 6061
rect 5944 5974 5978 5976
rect 5944 5938 5978 5940
rect 5944 5853 5978 5872
rect 6202 6042 6236 6061
rect 6202 5974 6236 5976
rect 6202 5938 6236 5940
rect 6202 5853 6236 5872
rect 6316 6003 6350 6037
rect 6316 5935 6350 5969
rect 6316 5867 6350 5901
rect 3508 5799 3542 5833
rect 3668 5785 3715 5819
rect 3751 5785 3785 5819
rect 3821 5785 3868 5819
rect 4442 5785 4489 5819
rect 4525 5785 4559 5819
rect 4595 5785 4642 5819
rect 4700 5785 4747 5819
rect 4783 5785 4817 5819
rect 4853 5785 4900 5819
rect 5474 5785 5521 5819
rect 5557 5785 5591 5819
rect 5627 5785 5674 5819
rect 5732 5785 5779 5819
rect 5815 5785 5849 5819
rect 5885 5785 5932 5819
rect 5990 5785 6037 5819
rect 6073 5785 6107 5819
rect 6143 5785 6190 5819
rect 6316 5799 6350 5833
rect 3508 5731 3542 5765
rect 6316 5731 6350 5765
rect 3508 5663 3542 5697
rect 3668 5677 3715 5711
rect 3751 5677 3785 5711
rect 3821 5677 3868 5711
rect 4442 5677 4489 5711
rect 4525 5677 4559 5711
rect 4595 5677 4642 5711
rect 4700 5677 4747 5711
rect 4783 5677 4817 5711
rect 4853 5677 4900 5711
rect 5474 5677 5521 5711
rect 5557 5677 5591 5711
rect 5627 5677 5674 5711
rect 5732 5677 5779 5711
rect 5815 5677 5849 5711
rect 5885 5677 5932 5711
rect 5990 5677 6037 5711
rect 6073 5677 6107 5711
rect 6143 5677 6190 5711
rect 6316 5663 6350 5697
rect 3508 5595 3542 5629
rect 3508 5527 3542 5561
rect 3508 5459 3542 5493
rect 3622 5624 3656 5643
rect 3622 5556 3656 5558
rect 3622 5520 3656 5522
rect 3622 5435 3656 5454
rect 3880 5624 3914 5643
rect 3880 5556 3914 5558
rect 3880 5520 3914 5522
rect 3880 5435 3914 5454
rect 4138 5624 4172 5643
rect 4138 5556 4172 5558
rect 4138 5520 4172 5522
rect 4138 5435 4172 5454
rect 4396 5624 4430 5643
rect 4396 5556 4430 5558
rect 4396 5520 4430 5522
rect 4396 5435 4430 5454
rect 4654 5624 4688 5643
rect 4654 5556 4688 5558
rect 4654 5520 4688 5522
rect 4654 5435 4688 5454
rect 4912 5624 4946 5643
rect 4912 5556 4946 5558
rect 4912 5520 4946 5522
rect 4912 5435 4946 5454
rect 5170 5624 5204 5643
rect 5170 5556 5204 5558
rect 5170 5520 5204 5522
rect 5170 5435 5204 5454
rect 5428 5624 5462 5643
rect 5428 5556 5462 5558
rect 5428 5520 5462 5522
rect 5428 5435 5462 5454
rect 5686 5624 5720 5643
rect 5686 5556 5720 5558
rect 5686 5520 5720 5522
rect 5686 5435 5720 5454
rect 5944 5624 5978 5643
rect 5944 5556 5978 5558
rect 5944 5520 5978 5522
rect 5944 5435 5978 5454
rect 6202 5624 6236 5643
rect 6202 5556 6236 5558
rect 6202 5520 6236 5522
rect 6202 5435 6236 5454
rect 6316 5595 6350 5629
rect 6316 5527 6350 5561
rect 6316 5459 6350 5493
rect 3508 5391 3542 5425
rect 3668 5367 3715 5401
rect 3751 5367 3785 5401
rect 3821 5367 3868 5401
rect 3926 5367 3973 5401
rect 4009 5367 4043 5401
rect 4079 5367 4126 5401
rect 4184 5367 4231 5401
rect 4267 5367 4301 5401
rect 4337 5367 4384 5401
rect 4958 5367 5005 5401
rect 5041 5367 5075 5401
rect 5111 5367 5158 5401
rect 5216 5367 5263 5401
rect 5299 5367 5333 5401
rect 5369 5367 5416 5401
rect 5990 5367 6037 5401
rect 6073 5367 6107 5401
rect 6143 5367 6190 5401
rect 6316 5391 6350 5425
rect 3508 5323 3542 5357
rect 6316 5323 6350 5357
rect 3508 5255 3542 5289
rect 3668 5259 3715 5293
rect 3751 5259 3785 5293
rect 3821 5259 3868 5293
rect 3926 5259 3973 5293
rect 4009 5259 4043 5293
rect 4079 5259 4126 5293
rect 4184 5259 4231 5293
rect 4267 5259 4301 5293
rect 4337 5259 4384 5293
rect 4958 5259 5005 5293
rect 5041 5259 5075 5293
rect 5111 5259 5158 5293
rect 5216 5259 5263 5293
rect 5299 5259 5333 5293
rect 5369 5259 5416 5293
rect 5990 5259 6037 5293
rect 6073 5259 6107 5293
rect 6143 5259 6190 5293
rect 6316 5255 6350 5289
rect 3508 5187 3542 5221
rect 3508 5119 3542 5153
rect 3508 5051 3542 5085
rect 3622 5206 3656 5225
rect 3622 5138 3656 5140
rect 3622 5102 3656 5104
rect 3622 5017 3656 5036
rect 3880 5206 3914 5225
rect 3880 5138 3914 5140
rect 3880 5102 3914 5104
rect 3880 5017 3914 5036
rect 4138 5206 4172 5225
rect 4138 5138 4172 5140
rect 4138 5102 4172 5104
rect 4138 5017 4172 5036
rect 4396 5206 4430 5225
rect 4396 5138 4430 5140
rect 4396 5102 4430 5104
rect 4396 5017 4430 5036
rect 4654 5206 4688 5225
rect 4654 5138 4688 5140
rect 4654 5102 4688 5104
rect 4654 5017 4688 5036
rect 4912 5206 4946 5225
rect 4912 5138 4946 5140
rect 4912 5102 4946 5104
rect 4912 5017 4946 5036
rect 5170 5206 5204 5225
rect 5170 5138 5204 5140
rect 5170 5102 5204 5104
rect 5170 5017 5204 5036
rect 5428 5206 5462 5225
rect 5428 5138 5462 5140
rect 5428 5102 5462 5104
rect 5428 5017 5462 5036
rect 5686 5206 5720 5225
rect 5686 5138 5720 5140
rect 5686 5102 5720 5104
rect 5686 5017 5720 5036
rect 5944 5206 5978 5225
rect 5944 5138 5978 5140
rect 5944 5102 5978 5104
rect 5944 5017 5978 5036
rect 6202 5206 6236 5225
rect 6202 5138 6236 5140
rect 6202 5102 6236 5104
rect 6202 5017 6236 5036
rect 6316 5187 6350 5221
rect 6316 5119 6350 5153
rect 6316 5051 6350 5085
rect 3508 4983 3542 5017
rect 3668 4949 3715 4983
rect 3751 4949 3785 4983
rect 3821 4949 3868 4983
rect 4442 4949 4489 4983
rect 4525 4949 4559 4983
rect 4595 4949 4642 4983
rect 4700 4949 4747 4983
rect 4783 4949 4817 4983
rect 4853 4949 4900 4983
rect 5474 4949 5521 4983
rect 5557 4949 5591 4983
rect 5627 4949 5674 4983
rect 5732 4949 5779 4983
rect 5815 4949 5849 4983
rect 5885 4949 5932 4983
rect 5990 4949 6037 4983
rect 6073 4949 6107 4983
rect 6143 4949 6190 4983
rect 3508 4915 3542 4949
rect 3508 4847 3542 4881
rect 6316 4915 6350 5017
rect 3668 4841 3715 4875
rect 3751 4841 3785 4875
rect 3821 4841 3868 4875
rect 4442 4841 4489 4875
rect 4525 4841 4559 4875
rect 4595 4841 4642 4875
rect 4700 4841 4747 4875
rect 4783 4841 4817 4875
rect 4853 4841 4900 4875
rect 5474 4841 5521 4875
rect 5557 4841 5591 4875
rect 5627 4841 5674 4875
rect 5732 4841 5779 4875
rect 5815 4841 5849 4875
rect 5885 4841 5932 4875
rect 5990 4841 6037 4875
rect 6073 4841 6107 4875
rect 6143 4841 6190 4875
rect 6316 4847 6350 4881
rect 3508 4779 3542 4813
rect 3508 4711 3542 4745
rect 3508 4643 3542 4677
rect 3508 4575 3542 4609
rect 3622 4788 3656 4807
rect 3622 4720 3656 4722
rect 3622 4684 3656 4686
rect 3622 4599 3656 4618
rect 3880 4788 3914 4807
rect 3880 4720 3914 4722
rect 3880 4684 3914 4686
rect 3880 4599 3914 4618
rect 4138 4788 4172 4807
rect 4138 4720 4172 4722
rect 4138 4684 4172 4686
rect 4138 4599 4172 4618
rect 4396 4788 4430 4807
rect 4396 4720 4430 4722
rect 4396 4684 4430 4686
rect 4396 4599 4430 4618
rect 4654 4788 4688 4807
rect 4654 4720 4688 4722
rect 4654 4684 4688 4686
rect 4654 4599 4688 4618
rect 4912 4788 4946 4807
rect 4912 4720 4946 4722
rect 4912 4684 4946 4686
rect 4912 4599 4946 4618
rect 5170 4788 5204 4807
rect 5170 4720 5204 4722
rect 5170 4684 5204 4686
rect 5170 4599 5204 4618
rect 5428 4788 5462 4807
rect 5428 4720 5462 4722
rect 5428 4684 5462 4686
rect 5428 4599 5462 4618
rect 5686 4788 5720 4807
rect 5686 4720 5720 4722
rect 5686 4684 5720 4686
rect 5686 4599 5720 4618
rect 5944 4788 5978 4807
rect 5944 4720 5978 4722
rect 5944 4684 5978 4686
rect 5944 4599 5978 4618
rect 6202 4788 6236 4807
rect 6202 4720 6236 4722
rect 6202 4684 6236 4686
rect 6202 4599 6236 4618
rect 6316 4779 6350 4813
rect 6316 4711 6350 4745
rect 6316 4643 6350 4677
rect 6316 4575 6350 4609
rect 3508 4507 3542 4541
rect 3668 4531 3715 4565
rect 3751 4531 3785 4565
rect 3821 4531 3868 4565
rect 3926 4531 3973 4565
rect 4009 4531 4043 4565
rect 4079 4531 4126 4565
rect 4184 4531 4231 4565
rect 4267 4531 4301 4565
rect 4337 4531 4384 4565
rect 4958 4531 5005 4565
rect 5041 4531 5075 4565
rect 5111 4531 5158 4565
rect 5216 4531 5263 4565
rect 5299 4531 5333 4565
rect 5369 4531 5416 4565
rect 5990 4531 6037 4565
rect 6073 4531 6107 4565
rect 6143 4531 6190 4565
rect 3508 4439 3542 4473
rect 6316 4507 6350 4541
rect 3668 4423 3715 4457
rect 3751 4423 3785 4457
rect 3821 4423 3868 4457
rect 3926 4423 3973 4457
rect 4009 4423 4043 4457
rect 4079 4423 4126 4457
rect 4184 4423 4231 4457
rect 4267 4423 4301 4457
rect 4337 4423 4384 4457
rect 4442 4423 4489 4457
rect 4525 4423 4559 4457
rect 4595 4423 4642 4457
rect 4700 4423 4747 4457
rect 4783 4423 4817 4457
rect 4853 4423 4900 4457
rect 4958 4423 5005 4457
rect 5041 4423 5075 4457
rect 5111 4423 5158 4457
rect 5216 4423 5263 4457
rect 5299 4423 5333 4457
rect 5369 4423 5416 4457
rect 5474 4423 5521 4457
rect 5557 4423 5591 4457
rect 5627 4423 5674 4457
rect 5732 4423 5779 4457
rect 5815 4423 5849 4457
rect 5885 4423 5932 4457
rect 5990 4423 6037 4457
rect 6073 4423 6107 4457
rect 6143 4423 6190 4457
rect 6316 4439 6350 4473
rect 3508 4371 3542 4405
rect 3508 4303 3542 4337
rect 3508 4235 3542 4269
rect 3508 4167 3542 4201
rect 3622 4370 3656 4389
rect 3622 4302 3656 4304
rect 3622 4266 3656 4268
rect 3622 4181 3656 4200
rect 3880 4370 3914 4389
rect 3880 4302 3914 4304
rect 3880 4266 3914 4268
rect 3880 4181 3914 4200
rect 4138 4370 4172 4389
rect 4138 4302 4172 4304
rect 4138 4266 4172 4268
rect 4138 4181 4172 4200
rect 4396 4370 4430 4389
rect 4396 4302 4430 4304
rect 4396 4266 4430 4268
rect 4396 4181 4430 4200
rect 4654 4370 4688 4389
rect 4654 4302 4688 4304
rect 4654 4266 4688 4268
rect 4654 4181 4688 4200
rect 4912 4370 4946 4389
rect 4912 4302 4946 4304
rect 4912 4266 4946 4268
rect 4912 4181 4946 4200
rect 5170 4370 5204 4389
rect 5170 4302 5204 4304
rect 5170 4266 5204 4268
rect 5170 4181 5204 4200
rect 5428 4370 5462 4389
rect 5428 4302 5462 4304
rect 5428 4266 5462 4268
rect 5428 4181 5462 4200
rect 5686 4370 5720 4389
rect 5686 4302 5720 4304
rect 5686 4266 5720 4268
rect 5686 4181 5720 4200
rect 5944 4370 5978 4389
rect 5944 4302 5978 4304
rect 5944 4266 5978 4268
rect 5944 4181 5978 4200
rect 6202 4370 6236 4389
rect 6202 4302 6236 4304
rect 6202 4266 6236 4268
rect 6202 4181 6236 4200
rect 6316 4371 6350 4405
rect 6316 4303 6350 4337
rect 6316 4238 6350 4269
rect 6316 4167 6350 4201
rect 3508 4045 3542 4133
rect 3668 4113 3715 4147
rect 3751 4113 3785 4147
rect 3821 4113 3868 4147
rect 5990 4113 6037 4147
rect 6073 4113 6107 4147
rect 6143 4113 6190 4147
rect 6316 4045 6350 4133
rect 3508 4011 3628 4045
rect 3662 4011 3696 4045
rect 3730 4011 3764 4045
rect 3798 4011 3832 4045
rect 3866 4011 3900 4045
rect 3934 4011 3968 4045
rect 4002 4011 4036 4045
rect 4070 4011 4104 4045
rect 4138 4011 4172 4045
rect 4206 4011 4240 4045
rect 4274 4011 4308 4045
rect 4342 4011 4376 4045
rect 4410 4011 4444 4045
rect 4478 4011 4512 4045
rect 4546 4011 4580 4045
rect 4614 4011 4648 4045
rect 4682 4011 4716 4045
rect 4750 4011 4784 4045
rect 4818 4011 4852 4045
rect 4886 4011 4920 4045
rect 4954 4011 4988 4045
rect 5022 4011 5056 4045
rect 5090 4011 5124 4045
rect 5158 4011 5192 4045
rect 5226 4011 5260 4045
rect 5294 4011 5328 4045
rect 5362 4011 5396 4045
rect 5430 4011 5464 4045
rect 5498 4011 5532 4045
rect 5566 4011 5600 4045
rect 5634 4011 5668 4045
rect 5702 4011 5736 4045
rect 5770 4011 5804 4045
rect 5838 4011 5872 4045
rect 5906 4011 5940 4045
rect 5974 4011 6008 4045
rect 6042 4011 6076 4045
rect 6110 4011 6144 4045
rect 6178 4011 6212 4045
rect 6246 4011 6350 4045
rect 8244 7040 8364 7074
rect 8398 7040 8432 7074
rect 8466 7040 8500 7074
rect 8534 7040 8568 7074
rect 8602 7040 8636 7074
rect 8670 7040 8704 7074
rect 8738 7040 8772 7074
rect 8806 7040 8840 7074
rect 8874 7040 8908 7074
rect 8942 7040 8976 7074
rect 9010 7040 9044 7074
rect 9078 7040 9112 7074
rect 9146 7040 9180 7074
rect 9214 7040 9248 7074
rect 9282 7040 9316 7074
rect 9350 7040 9384 7074
rect 9418 7040 9452 7074
rect 9486 7040 9520 7074
rect 9554 7040 9588 7074
rect 9622 7040 9656 7074
rect 9690 7040 9724 7074
rect 9758 7040 9792 7074
rect 9826 7040 9860 7074
rect 9894 7040 9928 7074
rect 9962 7040 10054 7074
rect 8244 6952 8278 7040
rect 8404 6938 8451 6972
rect 8487 6938 8521 6972
rect 8557 6938 8604 6972
rect 8662 6938 8709 6972
rect 8745 6938 8779 6972
rect 8815 6938 8862 6972
rect 8920 6938 8967 6972
rect 9003 6938 9037 6972
rect 9073 6938 9120 6972
rect 9178 6938 9225 6972
rect 9261 6938 9295 6972
rect 9331 6938 9378 6972
rect 9436 6938 9483 6972
rect 9519 6938 9553 6972
rect 9589 6938 9636 6972
rect 9694 6938 9741 6972
rect 9777 6938 9811 6972
rect 9847 6938 9894 6972
rect 10020 6952 10054 7040
rect 8244 6884 8278 6918
rect 8244 6816 8278 6850
rect 8244 6748 8278 6782
rect 8244 6680 8278 6714
rect 8358 6885 8392 6904
rect 8358 6817 8392 6819
rect 8358 6781 8392 6783
rect 8358 6696 8392 6715
rect 8616 6885 8650 6904
rect 8616 6817 8650 6819
rect 8616 6781 8650 6783
rect 8616 6696 8650 6715
rect 8874 6885 8908 6904
rect 8874 6817 8908 6819
rect 8874 6781 8908 6783
rect 8874 6696 8908 6715
rect 9132 6885 9166 6904
rect 9132 6817 9166 6819
rect 9132 6781 9166 6783
rect 9132 6696 9166 6715
rect 9390 6885 9424 6904
rect 9390 6817 9424 6819
rect 9390 6781 9424 6783
rect 9390 6696 9424 6715
rect 9648 6885 9682 6904
rect 9648 6817 9682 6819
rect 9648 6781 9682 6783
rect 9648 6696 9682 6715
rect 9906 6885 9940 6904
rect 9906 6817 9940 6819
rect 9906 6781 9940 6783
rect 9906 6696 9940 6715
rect 10020 6884 10054 6918
rect 10020 6816 10054 6850
rect 10020 6748 10054 6782
rect 10020 6680 10054 6714
rect 8244 6612 8278 6646
rect 8404 6628 8451 6662
rect 8487 6628 8521 6662
rect 8557 6628 8604 6662
rect 9694 6628 9741 6662
rect 9777 6628 9811 6662
rect 9847 6628 9894 6662
rect 8244 6544 8278 6578
rect 10020 6612 10054 6646
rect 8404 6520 8451 6554
rect 8487 6520 8521 6554
rect 8557 6520 8604 6554
rect 8662 6520 8709 6554
rect 8745 6520 8779 6554
rect 8815 6520 8862 6554
rect 8920 6520 8967 6554
rect 9003 6520 9037 6554
rect 9073 6520 9120 6554
rect 9178 6520 9225 6554
rect 9261 6520 9295 6554
rect 9331 6520 9378 6554
rect 9436 6520 9483 6554
rect 9519 6520 9553 6554
rect 9589 6520 9636 6554
rect 9694 6520 9741 6554
rect 9777 6520 9811 6554
rect 9847 6520 9894 6554
rect 10020 6544 10054 6578
rect 8244 6476 8278 6510
rect 8244 6408 8278 6442
rect 8244 6340 8278 6374
rect 8244 6272 8278 6306
rect 8358 6467 8392 6486
rect 8358 6399 8392 6401
rect 8358 6363 8392 6365
rect 8358 6278 8392 6297
rect 8616 6467 8650 6486
rect 8616 6399 8650 6401
rect 8616 6363 8650 6365
rect 8616 6278 8650 6297
rect 8874 6467 8908 6486
rect 8874 6399 8908 6401
rect 8874 6363 8908 6365
rect 8874 6278 8908 6297
rect 9132 6467 9166 6486
rect 9132 6399 9166 6401
rect 9132 6363 9166 6365
rect 9132 6278 9166 6297
rect 9390 6467 9424 6486
rect 9390 6399 9424 6401
rect 9390 6363 9424 6365
rect 9390 6278 9424 6297
rect 9648 6467 9682 6486
rect 9648 6399 9682 6401
rect 9648 6363 9682 6365
rect 9648 6278 9682 6297
rect 9906 6467 9940 6486
rect 9906 6399 9940 6401
rect 9906 6363 9940 6365
rect 9906 6278 9940 6297
rect 10020 6476 10054 6510
rect 10020 6408 10054 6442
rect 10020 6340 10054 6374
rect 10020 6272 10054 6306
rect 8244 6204 8278 6238
rect 8404 6210 8451 6244
rect 8487 6210 8521 6244
rect 8557 6210 8604 6244
rect 9694 6210 9741 6244
rect 9777 6210 9811 6244
rect 9847 6210 9894 6244
rect 8244 6136 8278 6170
rect 10020 6204 10054 6238
rect 8404 6102 8451 6136
rect 8487 6102 8521 6136
rect 8557 6102 8604 6136
rect 8662 6102 8709 6136
rect 8745 6102 8779 6136
rect 8815 6102 8862 6136
rect 8920 6102 8967 6136
rect 9003 6102 9037 6136
rect 9073 6102 9120 6136
rect 9178 6102 9225 6136
rect 9261 6102 9295 6136
rect 9331 6102 9378 6136
rect 9436 6102 9483 6136
rect 9519 6102 9553 6136
rect 9589 6102 9636 6136
rect 9694 6102 9741 6136
rect 9777 6102 9811 6136
rect 9847 6102 9894 6136
rect 8244 6068 8278 6102
rect 10020 6068 10054 6170
rect 8244 6000 8278 6034
rect 8244 5932 8278 5966
rect 8244 5864 8278 5898
rect 8358 6049 8392 6068
rect 8358 5981 8392 5983
rect 8358 5945 8392 5947
rect 8358 5860 8392 5879
rect 8616 6049 8650 6068
rect 8616 5981 8650 5983
rect 8616 5945 8650 5947
rect 8616 5860 8650 5879
rect 8874 6049 8908 6068
rect 8874 5981 8908 5983
rect 8874 5945 8908 5947
rect 8874 5860 8908 5879
rect 9132 6049 9166 6068
rect 9132 5981 9166 5983
rect 9132 5945 9166 5947
rect 9132 5860 9166 5879
rect 9390 6049 9424 6068
rect 9390 5981 9424 5983
rect 9390 5945 9424 5947
rect 9390 5860 9424 5879
rect 9648 6049 9682 6068
rect 9648 5981 9682 5983
rect 9648 5945 9682 5947
rect 9648 5860 9682 5879
rect 9906 6049 9940 6068
rect 9906 5981 9940 5983
rect 9906 5945 9940 5947
rect 9906 5860 9940 5879
rect 10020 6000 10054 6034
rect 10020 5932 10054 5966
rect 10020 5864 10054 5898
rect 8244 5796 8278 5830
rect 8404 5792 8451 5826
rect 8487 5792 8521 5826
rect 8557 5792 8604 5826
rect 9694 5792 9741 5826
rect 9777 5792 9811 5826
rect 9847 5792 9894 5826
rect 10020 5796 10054 5830
rect 8244 5728 8278 5762
rect 10020 5728 10054 5762
rect 8244 5660 8278 5694
rect 8404 5684 8451 5718
rect 8487 5684 8521 5718
rect 8557 5684 8604 5718
rect 8662 5684 8709 5718
rect 8745 5684 8779 5718
rect 8815 5684 8862 5718
rect 8920 5684 8967 5718
rect 9003 5684 9037 5718
rect 9073 5684 9120 5718
rect 9178 5684 9225 5718
rect 9261 5684 9295 5718
rect 9331 5684 9378 5718
rect 9436 5684 9483 5718
rect 9519 5684 9553 5718
rect 9589 5684 9636 5718
rect 9694 5684 9741 5718
rect 9777 5684 9811 5718
rect 9847 5684 9894 5718
rect 10020 5660 10054 5694
rect 8244 5592 8278 5626
rect 8244 5524 8278 5558
rect 8244 5456 8278 5490
rect 8358 5631 8392 5650
rect 8358 5563 8392 5565
rect 8358 5527 8392 5529
rect 8358 5442 8392 5461
rect 8616 5631 8650 5650
rect 8616 5563 8650 5565
rect 8616 5527 8650 5529
rect 8616 5442 8650 5461
rect 8874 5631 8908 5650
rect 8874 5563 8908 5565
rect 8874 5527 8908 5529
rect 8874 5442 8908 5461
rect 9132 5631 9166 5650
rect 9132 5563 9166 5565
rect 9132 5527 9166 5529
rect 9132 5442 9166 5461
rect 9390 5631 9424 5650
rect 9390 5563 9424 5565
rect 9390 5527 9424 5529
rect 9390 5442 9424 5461
rect 9648 5631 9682 5650
rect 9648 5563 9682 5565
rect 9648 5527 9682 5529
rect 9648 5442 9682 5461
rect 9906 5631 9940 5650
rect 9906 5563 9940 5565
rect 9906 5527 9940 5529
rect 9906 5442 9940 5461
rect 10020 5592 10054 5626
rect 10020 5524 10054 5558
rect 10020 5456 10054 5490
rect 8244 5388 8278 5422
rect 8404 5374 8451 5408
rect 8487 5374 8521 5408
rect 8557 5374 8604 5408
rect 9694 5374 9741 5408
rect 9777 5374 9811 5408
rect 9847 5374 9894 5408
rect 10020 5388 10054 5422
rect 8244 5320 8278 5354
rect 10020 5320 10054 5354
rect 8244 5252 8278 5286
rect 8404 5266 8451 5300
rect 8487 5266 8521 5300
rect 8557 5266 8604 5300
rect 8662 5266 8709 5300
rect 8745 5266 8779 5300
rect 8815 5266 8862 5300
rect 8920 5266 8967 5300
rect 9003 5266 9037 5300
rect 9073 5266 9120 5300
rect 9178 5266 9225 5300
rect 9261 5266 9295 5300
rect 9331 5266 9378 5300
rect 9436 5266 9483 5300
rect 9519 5266 9553 5300
rect 9589 5266 9636 5300
rect 9694 5266 9741 5300
rect 9777 5266 9811 5300
rect 9847 5266 9894 5300
rect 10020 5252 10054 5286
rect 8244 5184 8278 5218
rect 8244 5116 8278 5150
rect 8244 5048 8278 5082
rect 8358 5213 8392 5232
rect 8358 5145 8392 5147
rect 8358 5109 8392 5111
rect 8358 5024 8392 5043
rect 8616 5213 8650 5232
rect 8616 5145 8650 5147
rect 8616 5109 8650 5111
rect 8616 5024 8650 5043
rect 8874 5213 8908 5232
rect 8874 5145 8908 5147
rect 8874 5109 8908 5111
rect 8874 5024 8908 5043
rect 9132 5213 9166 5232
rect 9132 5145 9166 5147
rect 9132 5109 9166 5111
rect 9132 5024 9166 5043
rect 9390 5213 9424 5232
rect 9390 5145 9424 5147
rect 9390 5109 9424 5111
rect 9390 5024 9424 5043
rect 9648 5213 9682 5232
rect 9648 5145 9682 5147
rect 9648 5109 9682 5111
rect 9648 5024 9682 5043
rect 9906 5213 9940 5232
rect 9906 5145 9940 5147
rect 9906 5109 9940 5111
rect 9906 5024 9940 5043
rect 10020 5184 10054 5218
rect 10020 5116 10054 5150
rect 10020 5048 10054 5082
rect 8244 4980 8278 5014
rect 8404 4956 8451 4990
rect 8487 4956 8521 4990
rect 8557 4956 8604 4990
rect 9694 4956 9741 4990
rect 9777 4956 9811 4990
rect 9847 4956 9894 4990
rect 10020 4980 10054 5014
rect 8244 4912 8278 4946
rect 10020 4912 10054 4946
rect 8244 4844 8278 4878
rect 8404 4848 8451 4882
rect 8487 4848 8521 4882
rect 8557 4848 8604 4882
rect 8662 4848 8709 4882
rect 8745 4848 8779 4882
rect 8815 4848 8862 4882
rect 8920 4848 8967 4882
rect 9003 4848 9037 4882
rect 9073 4848 9120 4882
rect 9178 4848 9225 4882
rect 9261 4848 9295 4882
rect 9331 4848 9378 4882
rect 9436 4848 9483 4882
rect 9519 4848 9553 4882
rect 9589 4848 9636 4882
rect 9694 4848 9741 4882
rect 9777 4848 9811 4882
rect 9847 4848 9894 4882
rect 10020 4844 10054 4878
rect 8244 4776 8278 4810
rect 8244 4708 8278 4742
rect 8244 4640 8278 4674
rect 8358 4795 8392 4814
rect 8358 4727 8392 4729
rect 8358 4691 8392 4693
rect 8358 4606 8392 4625
rect 8616 4795 8650 4814
rect 8616 4727 8650 4729
rect 8616 4691 8650 4693
rect 8616 4606 8650 4625
rect 8874 4795 8908 4814
rect 8874 4727 8908 4729
rect 8874 4691 8908 4693
rect 8874 4606 8908 4625
rect 9132 4795 9166 4814
rect 9132 4727 9166 4729
rect 9132 4691 9166 4693
rect 9132 4606 9166 4625
rect 9390 4795 9424 4814
rect 9390 4727 9424 4729
rect 9390 4691 9424 4693
rect 9390 4606 9424 4625
rect 9648 4795 9682 4814
rect 9648 4727 9682 4729
rect 9648 4691 9682 4693
rect 9648 4606 9682 4625
rect 9906 4795 9940 4814
rect 9906 4727 9940 4729
rect 9906 4691 9940 4693
rect 9906 4606 9940 4625
rect 10020 4776 10054 4810
rect 10020 4708 10054 4742
rect 10020 4640 10054 4674
rect 8244 4572 8278 4606
rect 8404 4538 8451 4572
rect 8487 4538 8521 4572
rect 8557 4538 8604 4572
rect 9694 4538 9741 4572
rect 9777 4538 9811 4572
rect 9847 4538 9894 4572
rect 8244 4504 8278 4538
rect 8244 4436 8278 4470
rect 10020 4504 10054 4606
rect 8404 4430 8451 4464
rect 8487 4430 8521 4464
rect 8557 4430 8604 4464
rect 8662 4430 8709 4464
rect 8745 4430 8779 4464
rect 8815 4430 8862 4464
rect 8920 4430 8967 4464
rect 9003 4430 9037 4464
rect 9073 4430 9120 4464
rect 9178 4430 9225 4464
rect 9261 4430 9295 4464
rect 9331 4430 9378 4464
rect 9436 4430 9483 4464
rect 9519 4430 9553 4464
rect 9589 4430 9636 4464
rect 9694 4430 9741 4464
rect 9777 4430 9811 4464
rect 9847 4430 9894 4464
rect 10020 4436 10054 4470
rect 8244 4368 8278 4402
rect 8244 4300 8278 4334
rect 8244 4232 8278 4266
rect 8244 4164 8278 4198
rect 8358 4377 8392 4396
rect 8358 4309 8392 4311
rect 8358 4273 8392 4275
rect 8358 4188 8392 4207
rect 8616 4377 8650 4396
rect 8616 4309 8650 4311
rect 8616 4273 8650 4275
rect 8616 4188 8650 4207
rect 8874 4377 8908 4396
rect 8874 4309 8908 4311
rect 8874 4273 8908 4275
rect 8874 4188 8908 4207
rect 9132 4377 9166 4396
rect 9132 4309 9166 4311
rect 9132 4273 9166 4275
rect 9132 4188 9166 4207
rect 9390 4377 9424 4396
rect 9390 4309 9424 4311
rect 9390 4273 9424 4275
rect 9390 4188 9424 4207
rect 9648 4377 9682 4396
rect 9648 4309 9682 4311
rect 9648 4273 9682 4275
rect 9648 4188 9682 4207
rect 9906 4377 9940 4396
rect 9906 4309 9940 4311
rect 9906 4273 9940 4275
rect 9906 4188 9940 4207
rect 10020 4368 10054 4402
rect 10020 4300 10054 4334
rect 10020 4232 10054 4266
rect 10020 4164 10054 4198
rect 8244 4052 8278 4130
rect 8404 4120 8451 4154
rect 8487 4120 8521 4154
rect 8557 4120 8604 4154
rect 9694 4120 9741 4154
rect 9777 4120 9811 4154
rect 9847 4120 9894 4154
rect 10020 4052 10054 4130
rect 8244 4018 8364 4052
rect 8398 4018 8432 4052
rect 8466 4018 8500 4052
rect 8534 4018 8568 4052
rect 8602 4018 8636 4052
rect 8670 4018 8704 4052
rect 8738 4018 8772 4052
rect 8806 4018 8840 4052
rect 8874 4018 8908 4052
rect 8942 4018 8976 4052
rect 9010 4018 9044 4052
rect 9078 4018 9112 4052
rect 9146 4018 9180 4052
rect 9214 4018 9248 4052
rect 9282 4018 9316 4052
rect 9350 4018 9384 4052
rect 9418 4018 9452 4052
rect 9486 4018 9520 4052
rect 9554 4018 9588 4052
rect 9622 4018 9656 4052
rect 9690 4018 9724 4052
rect 9758 4018 9792 4052
rect 9826 4018 9860 4052
rect 9894 4018 9906 4052
rect 9940 4018 10054 4052
rect 1518 3990 1552 4007
rect -2322 3848 -2288 3956
rect -2162 3916 -2115 3950
rect -2079 3916 -2045 3950
rect -2009 3916 -1962 3950
rect 1192 3916 1239 3950
rect 1275 3916 1309 3950
rect 1345 3916 1392 3950
rect 1518 3848 1552 3956
rect -2322 3814 -2202 3848
rect -2168 3814 -2134 3848
rect -2100 3814 -2066 3848
rect -2032 3814 -1998 3848
rect -1964 3814 -1930 3848
rect -1896 3814 -1862 3848
rect -1828 3814 -1794 3848
rect -1760 3814 -1726 3848
rect -1692 3814 -1658 3848
rect -1624 3814 -1590 3848
rect -1556 3814 -1522 3848
rect -1488 3814 -1454 3848
rect -1420 3814 -1386 3848
rect -1352 3814 -1318 3848
rect -1284 3814 -1250 3848
rect -1216 3814 -1182 3848
rect -1148 3814 -1114 3848
rect -1080 3814 -1046 3848
rect -1012 3814 -978 3848
rect -944 3814 -910 3848
rect -876 3814 -842 3848
rect -808 3814 -774 3848
rect -740 3814 -706 3848
rect -672 3814 -638 3848
rect -604 3814 -570 3848
rect -536 3814 -502 3848
rect -468 3814 -434 3848
rect -400 3814 -366 3848
rect -332 3814 -298 3848
rect -264 3814 -230 3848
rect -196 3814 -162 3848
rect -128 3814 -94 3848
rect -60 3814 -26 3848
rect 8 3814 42 3848
rect 76 3814 110 3848
rect 144 3814 178 3848
rect 212 3814 246 3848
rect 280 3814 314 3848
rect 348 3814 382 3848
rect 416 3814 450 3848
rect 484 3814 518 3848
rect 552 3814 586 3848
rect 620 3814 654 3848
rect 688 3814 722 3848
rect 756 3814 790 3848
rect 824 3814 858 3848
rect 892 3814 926 3848
rect 960 3814 994 3848
rect 1028 3814 1062 3848
rect 1096 3814 1130 3848
rect 1164 3814 1198 3848
rect 1232 3814 1266 3848
rect 1300 3814 1334 3848
rect 1368 3814 1402 3848
rect 1436 3814 1552 3848
<< viali >>
rect 8299 10947 8307 10981
rect 8307 10947 8333 10981
rect 3176 10737 3178 10771
rect 3178 10737 3210 10771
rect 3248 10737 3280 10771
rect 3280 10737 3282 10771
rect 3434 10737 3436 10771
rect 3436 10737 3468 10771
rect 3506 10737 3538 10771
rect 3538 10737 3540 10771
rect 3692 10737 3694 10771
rect 3694 10737 3726 10771
rect 3764 10737 3796 10771
rect 3796 10737 3798 10771
rect 4466 10737 4468 10771
rect 4468 10737 4500 10771
rect 4538 10737 4570 10771
rect 4570 10737 4572 10771
rect 4724 10737 4726 10771
rect 4726 10737 4758 10771
rect 4796 10737 4828 10771
rect 4828 10737 4830 10771
rect 4982 10737 4984 10771
rect 4984 10737 5016 10771
rect 5054 10737 5086 10771
rect 5086 10737 5088 10771
rect -1239 10629 -1233 10663
rect -1233 10629 -1205 10663
rect -1146 10527 -1144 10561
rect -1144 10527 -1112 10561
rect -1074 10527 -1042 10561
rect -1042 10527 -1040 10561
rect 144 10527 146 10561
rect 146 10527 178 10561
rect 216 10527 248 10561
rect 248 10527 250 10561
rect -1239 10431 -1205 10433
rect -1239 10399 -1205 10431
rect -1239 10329 -1205 10361
rect -1239 10327 -1205 10329
rect -981 10431 -947 10433
rect -981 10399 -947 10431
rect -981 10329 -947 10361
rect -981 10327 -947 10329
rect -723 10431 -689 10433
rect -723 10399 -689 10431
rect -723 10329 -689 10361
rect -723 10327 -689 10329
rect -465 10431 -431 10433
rect -465 10399 -431 10431
rect -465 10329 -431 10361
rect -465 10327 -431 10329
rect -207 10431 -173 10433
rect -207 10399 -173 10431
rect -207 10329 -173 10361
rect -207 10327 -173 10329
rect 51 10431 85 10433
rect 51 10399 85 10431
rect 51 10329 85 10361
rect 51 10327 85 10329
rect 309 10431 343 10433
rect 309 10399 343 10431
rect 309 10329 343 10361
rect 309 10327 343 10329
rect -1146 10199 -1144 10233
rect -1144 10199 -1112 10233
rect -1074 10199 -1042 10233
rect -1042 10199 -1040 10233
rect -888 10199 -886 10233
rect -886 10199 -854 10233
rect -816 10199 -784 10233
rect -784 10199 -782 10233
rect -630 10199 -628 10233
rect -628 10199 -596 10233
rect -558 10199 -526 10233
rect -526 10199 -524 10233
rect -372 10199 -370 10233
rect -370 10199 -338 10233
rect -300 10199 -268 10233
rect -268 10199 -266 10233
rect -114 10199 -112 10233
rect -112 10199 -80 10233
rect -42 10199 -10 10233
rect -10 10199 -8 10233
rect 144 10199 146 10233
rect 146 10199 178 10233
rect 216 10199 248 10233
rect 248 10199 250 10233
rect -1146 10091 -1144 10125
rect -1144 10091 -1112 10125
rect -1074 10091 -1042 10125
rect -1042 10091 -1040 10125
rect -888 10091 -886 10125
rect -886 10091 -854 10125
rect -816 10091 -784 10125
rect -784 10091 -782 10125
rect -630 10091 -628 10125
rect -628 10091 -596 10125
rect -558 10091 -526 10125
rect -526 10091 -524 10125
rect -372 10091 -370 10125
rect -370 10091 -338 10125
rect -300 10091 -268 10125
rect -268 10091 -266 10125
rect -114 10091 -112 10125
rect -112 10091 -80 10125
rect -42 10091 -10 10125
rect -10 10091 -8 10125
rect 144 10091 146 10125
rect 146 10091 178 10125
rect 216 10091 248 10125
rect 248 10091 250 10125
rect -1239 9995 -1205 9997
rect -1239 9963 -1205 9995
rect -1239 9893 -1205 9925
rect -1239 9891 -1205 9893
rect -981 9995 -947 9997
rect -981 9963 -947 9995
rect -981 9893 -947 9925
rect -981 9891 -947 9893
rect -723 9995 -689 9997
rect -723 9963 -689 9995
rect -723 9893 -689 9925
rect -723 9891 -689 9893
rect -465 9995 -431 9997
rect -465 9963 -431 9995
rect -465 9893 -431 9925
rect -465 9891 -431 9893
rect -207 9995 -173 9997
rect -207 9963 -173 9995
rect -207 9893 -173 9925
rect -207 9891 -173 9893
rect 51 9995 85 9997
rect 51 9963 85 9995
rect 51 9893 85 9925
rect 51 9891 85 9893
rect 309 9995 343 9997
rect 309 9963 343 9995
rect 309 9893 343 9925
rect 309 9891 343 9893
rect -1146 9763 -1144 9797
rect -1144 9763 -1112 9797
rect -1074 9763 -1042 9797
rect -1042 9763 -1040 9797
rect 144 9763 146 9797
rect 146 9763 178 9797
rect 216 9763 248 9797
rect 248 9763 250 9797
rect -1146 9655 -1144 9689
rect -1144 9655 -1112 9689
rect -1074 9655 -1042 9689
rect -1042 9655 -1040 9689
rect 144 9655 146 9689
rect 146 9655 178 9689
rect 216 9655 248 9689
rect 248 9655 250 9689
rect -1239 9559 -1205 9561
rect -1239 9527 -1205 9559
rect -1239 9457 -1205 9489
rect -1239 9455 -1205 9457
rect -981 9559 -947 9561
rect -981 9527 -947 9559
rect -981 9457 -947 9489
rect -981 9455 -947 9457
rect -723 9559 -689 9561
rect -723 9527 -689 9559
rect -723 9457 -689 9489
rect -723 9455 -689 9457
rect -465 9559 -431 9561
rect -465 9527 -431 9559
rect -465 9457 -431 9489
rect -465 9455 -431 9457
rect -207 9559 -173 9561
rect -207 9527 -173 9559
rect -207 9457 -173 9489
rect -207 9455 -173 9457
rect 51 9559 85 9561
rect 51 9527 85 9559
rect 51 9457 85 9489
rect 51 9455 85 9457
rect 309 9559 343 9561
rect 309 9527 343 9559
rect 309 9457 343 9489
rect 309 9455 343 9457
rect -1146 9327 -1144 9361
rect -1144 9327 -1112 9361
rect -1074 9327 -1042 9361
rect -1042 9327 -1040 9361
rect -888 9327 -886 9361
rect -886 9327 -854 9361
rect -816 9327 -784 9361
rect -784 9327 -782 9361
rect -630 9327 -628 9361
rect -628 9327 -596 9361
rect -558 9327 -526 9361
rect -526 9327 -524 9361
rect -372 9327 -370 9361
rect -370 9327 -338 9361
rect -300 9327 -268 9361
rect -268 9327 -266 9361
rect -114 9327 -112 9361
rect -112 9327 -80 9361
rect -42 9327 -10 9361
rect -10 9327 -8 9361
rect 144 9327 146 9361
rect 146 9327 178 9361
rect 216 9327 248 9361
rect 248 9327 250 9361
rect -1146 9219 -1144 9253
rect -1144 9219 -1112 9253
rect -1074 9219 -1042 9253
rect -1042 9219 -1040 9253
rect -888 9219 -886 9253
rect -886 9219 -854 9253
rect -816 9219 -784 9253
rect -784 9219 -782 9253
rect -630 9219 -628 9253
rect -628 9219 -596 9253
rect -558 9219 -526 9253
rect -526 9219 -524 9253
rect -372 9219 -370 9253
rect -370 9219 -338 9253
rect -300 9219 -268 9253
rect -268 9219 -266 9253
rect -114 9219 -112 9253
rect -112 9219 -80 9253
rect -42 9219 -10 9253
rect -10 9219 -8 9253
rect 144 9219 146 9253
rect 146 9219 178 9253
rect 216 9219 248 9253
rect 248 9219 250 9253
rect -1239 9123 -1205 9125
rect -1239 9091 -1205 9123
rect -1239 9021 -1205 9053
rect -1239 9019 -1205 9021
rect -981 9123 -947 9125
rect -981 9091 -947 9123
rect -981 9021 -947 9053
rect -981 9019 -947 9021
rect -723 9123 -689 9125
rect -723 9091 -689 9123
rect -723 9021 -689 9053
rect -723 9019 -689 9021
rect -465 9123 -431 9125
rect -465 9091 -431 9123
rect -465 9021 -431 9053
rect -465 9019 -431 9021
rect -207 9123 -173 9125
rect -207 9091 -173 9123
rect -207 9021 -173 9053
rect -207 9019 -173 9021
rect 51 9123 85 9125
rect 51 9091 85 9123
rect 51 9021 85 9053
rect 51 9019 85 9021
rect 309 9123 343 9125
rect 309 9091 343 9123
rect 309 9021 343 9053
rect 309 9019 343 9021
rect -1146 8891 -1144 8925
rect -1144 8891 -1112 8925
rect -1074 8891 -1042 8925
rect -1042 8891 -1040 8925
rect 144 8891 146 8925
rect 146 8891 178 8925
rect 216 8891 248 8925
rect 248 8891 250 8925
rect 3083 10650 3117 10652
rect 3083 10618 3117 10650
rect 3083 10548 3117 10580
rect 3083 10546 3117 10548
rect 3341 10650 3375 10652
rect 3341 10618 3375 10650
rect 3341 10548 3375 10580
rect 3341 10546 3375 10548
rect 3599 10650 3633 10652
rect 3599 10618 3633 10650
rect 3599 10548 3633 10580
rect 3599 10546 3633 10548
rect 3857 10650 3891 10652
rect 3857 10618 3891 10650
rect 3857 10548 3891 10580
rect 3857 10546 3891 10548
rect 4115 10650 4149 10652
rect 4115 10618 4149 10650
rect 4115 10548 4149 10580
rect 4115 10546 4149 10548
rect 4373 10650 4407 10652
rect 4373 10618 4407 10650
rect 4373 10548 4407 10580
rect 4373 10546 4407 10548
rect 4631 10650 4665 10652
rect 4631 10618 4665 10650
rect 4631 10548 4665 10580
rect 4631 10546 4665 10548
rect 4889 10650 4923 10652
rect 4889 10618 4923 10650
rect 4889 10548 4923 10580
rect 4889 10546 4923 10548
rect 5147 10650 5181 10652
rect 5147 10618 5181 10650
rect 5147 10548 5181 10580
rect 5147 10546 5181 10548
rect 3176 10427 3178 10461
rect 3178 10427 3210 10461
rect 3248 10427 3280 10461
rect 3280 10427 3282 10461
rect 3950 10427 3952 10461
rect 3952 10427 3984 10461
rect 4022 10427 4054 10461
rect 4054 10427 4056 10461
rect 4208 10427 4210 10461
rect 4210 10427 4242 10461
rect 4280 10427 4312 10461
rect 4312 10427 4314 10461
rect 4982 10424 4984 10458
rect 4984 10424 5016 10458
rect 5054 10424 5086 10458
rect 5086 10424 5088 10458
rect 3176 10319 3178 10353
rect 3178 10319 3210 10353
rect 3248 10319 3280 10353
rect 3280 10319 3282 10353
rect 3950 10319 3952 10353
rect 3952 10319 3984 10353
rect 4022 10319 4054 10353
rect 4054 10319 4056 10353
rect 4208 10319 4210 10353
rect 4210 10319 4242 10353
rect 4280 10319 4312 10353
rect 4312 10319 4314 10353
rect 4982 10319 4984 10353
rect 4984 10319 5016 10353
rect 5054 10319 5086 10353
rect 5086 10319 5088 10353
rect 3083 10232 3117 10234
rect 3083 10200 3117 10232
rect 3083 10130 3117 10162
rect 3083 10128 3117 10130
rect 3341 10232 3375 10234
rect 3341 10200 3375 10232
rect 3341 10130 3375 10162
rect 3341 10128 3375 10130
rect 3599 10232 3633 10234
rect 3599 10200 3633 10232
rect 3599 10130 3633 10162
rect 3599 10128 3633 10130
rect 3857 10232 3891 10234
rect 3857 10200 3891 10232
rect 3857 10130 3891 10162
rect 3857 10128 3891 10130
rect 4115 10232 4149 10234
rect 4115 10200 4149 10232
rect 4115 10130 4149 10162
rect 4115 10128 4149 10130
rect 4373 10232 4407 10234
rect 4373 10200 4407 10232
rect 4373 10130 4407 10162
rect 4373 10128 4407 10130
rect 4631 10232 4665 10234
rect 4631 10200 4665 10232
rect 4631 10130 4665 10162
rect 4631 10128 4665 10130
rect 4889 10232 4923 10234
rect 4889 10200 4923 10232
rect 4889 10130 4923 10162
rect 4889 10128 4923 10130
rect 5147 10232 5181 10234
rect 5147 10200 5181 10232
rect 5147 10130 5181 10162
rect 5147 10128 5181 10130
rect 3176 10009 3178 10043
rect 3178 10009 3210 10043
rect 3248 10009 3280 10043
rect 3280 10009 3282 10043
rect 3434 10009 3436 10043
rect 3436 10009 3468 10043
rect 3506 10009 3538 10043
rect 3538 10009 3540 10043
rect 3692 10009 3694 10043
rect 3694 10009 3726 10043
rect 3764 10009 3796 10043
rect 3796 10009 3798 10043
rect 4466 10009 4468 10043
rect 4468 10009 4500 10043
rect 4538 10009 4570 10043
rect 4570 10009 4572 10043
rect 4724 10009 4726 10043
rect 4726 10009 4758 10043
rect 4796 10009 4828 10043
rect 4828 10009 4830 10043
rect 4982 10009 4984 10043
rect 4984 10009 5016 10043
rect 5054 10009 5086 10043
rect 5086 10009 5088 10043
rect 3176 9901 3178 9935
rect 3178 9901 3210 9935
rect 3248 9901 3280 9935
rect 3280 9901 3282 9935
rect 3434 9901 3436 9935
rect 3436 9901 3468 9935
rect 3506 9901 3538 9935
rect 3538 9901 3540 9935
rect 3692 9901 3694 9935
rect 3694 9901 3726 9935
rect 3764 9901 3796 9935
rect 3796 9901 3798 9935
rect 4466 9901 4468 9935
rect 4468 9901 4500 9935
rect 4538 9901 4570 9935
rect 4570 9901 4572 9935
rect 4724 9901 4726 9935
rect 4726 9901 4758 9935
rect 4796 9901 4828 9935
rect 4828 9901 4830 9935
rect 4982 9901 4984 9935
rect 4984 9901 5016 9935
rect 5054 9901 5086 9935
rect 5086 9901 5088 9935
rect 3083 9814 3117 9816
rect 3083 9782 3117 9814
rect 3083 9712 3117 9744
rect 3083 9710 3117 9712
rect 3341 9814 3375 9816
rect 3341 9782 3375 9814
rect 3341 9712 3375 9744
rect 3341 9710 3375 9712
rect 3599 9814 3633 9816
rect 3599 9782 3633 9814
rect 3599 9712 3633 9744
rect 3599 9710 3633 9712
rect 3857 9814 3891 9816
rect 3857 9782 3891 9814
rect 3857 9712 3891 9744
rect 3857 9710 3891 9712
rect 4115 9814 4149 9816
rect 4115 9782 4149 9814
rect 4115 9712 4149 9744
rect 4115 9710 4149 9712
rect 4373 9814 4407 9816
rect 4373 9782 4407 9814
rect 4373 9712 4407 9744
rect 4373 9710 4407 9712
rect 4631 9814 4665 9816
rect 4631 9782 4665 9814
rect 4631 9712 4665 9744
rect 4631 9710 4665 9712
rect 4889 9814 4923 9816
rect 4889 9782 4923 9814
rect 4889 9712 4923 9744
rect 4889 9710 4923 9712
rect 5147 9814 5181 9816
rect 5147 9782 5181 9814
rect 5147 9712 5181 9744
rect 5147 9710 5181 9712
rect 3176 9591 3178 9625
rect 3178 9591 3210 9625
rect 3248 9591 3280 9625
rect 3280 9591 3282 9625
rect 3950 9591 3952 9625
rect 3952 9591 3984 9625
rect 4022 9591 4054 9625
rect 4054 9591 4056 9625
rect 4208 9591 4210 9625
rect 4210 9591 4242 9625
rect 4280 9591 4312 9625
rect 4312 9591 4314 9625
rect 4982 9588 4984 9622
rect 4984 9588 5016 9622
rect 5054 9588 5086 9622
rect 5086 9588 5088 9622
rect 3176 9483 3178 9517
rect 3178 9483 3210 9517
rect 3248 9483 3280 9517
rect 3280 9483 3282 9517
rect 3950 9483 3952 9517
rect 3952 9483 3984 9517
rect 4022 9483 4054 9517
rect 4054 9483 4056 9517
rect 4208 9483 4210 9517
rect 4210 9483 4242 9517
rect 4280 9483 4312 9517
rect 4312 9483 4314 9517
rect 4982 9483 4984 9517
rect 4984 9483 5016 9517
rect 5054 9483 5086 9517
rect 5086 9483 5088 9517
rect 3083 9396 3117 9398
rect 3083 9364 3117 9396
rect 3083 9294 3117 9326
rect 3083 9292 3117 9294
rect 3341 9396 3375 9398
rect 3341 9364 3375 9396
rect 3341 9294 3375 9326
rect 3341 9292 3375 9294
rect 3599 9396 3633 9398
rect 3599 9364 3633 9396
rect 3599 9294 3633 9326
rect 3599 9292 3633 9294
rect 3857 9396 3891 9398
rect 3857 9364 3891 9396
rect 3857 9294 3891 9326
rect 3857 9292 3891 9294
rect 4115 9396 4149 9398
rect 4115 9364 4149 9396
rect 4115 9294 4149 9326
rect 4115 9292 4149 9294
rect 4373 9396 4407 9398
rect 4373 9364 4407 9396
rect 4373 9294 4407 9326
rect 4373 9292 4407 9294
rect 4631 9396 4665 9398
rect 4631 9364 4665 9396
rect 4631 9294 4665 9326
rect 4631 9292 4665 9294
rect 4889 9396 4923 9398
rect 4889 9364 4923 9396
rect 4889 9294 4923 9326
rect 4889 9292 4923 9294
rect 5147 9396 5181 9398
rect 5147 9364 5181 9396
rect 5147 9294 5181 9326
rect 5147 9292 5181 9294
rect 3176 9173 3178 9207
rect 3178 9173 3210 9207
rect 3248 9173 3280 9207
rect 3280 9173 3282 9207
rect 3434 9173 3436 9207
rect 3436 9173 3468 9207
rect 3506 9173 3538 9207
rect 3538 9173 3540 9207
rect 3692 9173 3694 9207
rect 3694 9173 3726 9207
rect 3764 9173 3796 9207
rect 3796 9173 3798 9207
rect 4466 9173 4468 9207
rect 4468 9173 4500 9207
rect 4538 9173 4570 9207
rect 4570 9173 4572 9207
rect 4724 9173 4726 9207
rect 4726 9173 4758 9207
rect 4796 9173 4828 9207
rect 4828 9173 4830 9207
rect 4982 9170 4984 9204
rect 4984 9170 5016 9204
rect 5054 9170 5086 9204
rect 5086 9170 5088 9204
rect 3176 9061 3178 9095
rect 3178 9061 3210 9095
rect 3248 9061 3280 9095
rect 3280 9061 3282 9095
rect 3434 9061 3436 9095
rect 3436 9061 3468 9095
rect 3506 9061 3538 9095
rect 3538 9061 3540 9095
rect 3692 9061 3694 9095
rect 3694 9061 3726 9095
rect 3764 9061 3796 9095
rect 3796 9061 3798 9095
rect 4466 9061 4468 9095
rect 4468 9061 4500 9095
rect 4538 9061 4570 9095
rect 4570 9061 4572 9095
rect 4724 9061 4726 9095
rect 4726 9061 4758 9095
rect 4796 9061 4828 9095
rect 4828 9061 4830 9095
rect 4982 9061 4984 9095
rect 4984 9061 5016 9095
rect 5054 9061 5086 9095
rect 5086 9061 5088 9095
rect 3083 8974 3117 8976
rect 3083 8942 3117 8974
rect 3083 8872 3117 8904
rect 3083 8870 3117 8872
rect 3341 8974 3375 8976
rect 3341 8942 3375 8974
rect 3341 8872 3375 8904
rect 3341 8870 3375 8872
rect 3599 8974 3633 8976
rect 3599 8942 3633 8974
rect 3599 8872 3633 8904
rect 3599 8870 3633 8872
rect 3857 8974 3891 8976
rect 3857 8942 3891 8974
rect 3857 8872 3891 8904
rect 3857 8870 3891 8872
rect 4115 8974 4149 8976
rect 4115 8942 4149 8974
rect 4115 8872 4149 8904
rect 4115 8870 4149 8872
rect 4373 8974 4407 8976
rect 4373 8942 4407 8974
rect 4373 8872 4407 8904
rect 4373 8870 4407 8872
rect 4631 8974 4665 8976
rect 4631 8942 4665 8974
rect 4631 8872 4665 8904
rect 4631 8870 4665 8872
rect 4889 8974 4923 8976
rect 4889 8942 4923 8974
rect 4889 8872 4923 8904
rect 4889 8870 4923 8872
rect 5147 8974 5181 8976
rect 5147 8942 5181 8974
rect 5147 8872 5181 8904
rect 5147 8870 5181 8872
rect 3176 8751 3178 8785
rect 3178 8751 3210 8785
rect 3248 8751 3280 8785
rect 3280 8751 3282 8785
rect 3950 8751 3952 8785
rect 3952 8751 3984 8785
rect 4022 8751 4054 8785
rect 4054 8751 4056 8785
rect 4208 8751 4210 8785
rect 4210 8751 4242 8785
rect 4280 8751 4312 8785
rect 4312 8751 4314 8785
rect 4982 8748 4984 8782
rect 4984 8748 5016 8782
rect 5054 8748 5086 8782
rect 5086 8748 5088 8782
rect 3176 8639 3178 8673
rect 3178 8639 3210 8673
rect 3248 8639 3280 8673
rect 3280 8639 3282 8673
rect 3950 8639 3952 8673
rect 3952 8639 3984 8673
rect 4022 8639 4054 8673
rect 4054 8639 4056 8673
rect 4208 8639 4210 8673
rect 4210 8639 4242 8673
rect 4280 8639 4312 8673
rect 4312 8639 4314 8673
rect 4982 8639 4984 8673
rect 4984 8639 5016 8673
rect 5054 8639 5086 8673
rect 5086 8639 5088 8673
rect 3083 8552 3117 8554
rect 3083 8520 3117 8552
rect 3083 8450 3117 8482
rect 3083 8448 3117 8450
rect 3341 8552 3375 8554
rect 3341 8520 3375 8552
rect 3341 8450 3375 8482
rect 3341 8448 3375 8450
rect 3599 8552 3633 8554
rect 3599 8520 3633 8552
rect 3599 8450 3633 8482
rect 3599 8448 3633 8450
rect 3857 8552 3891 8554
rect 3857 8520 3891 8552
rect 3857 8450 3891 8482
rect 3857 8448 3891 8450
rect 4115 8552 4149 8554
rect 4115 8520 4149 8552
rect 4115 8450 4149 8482
rect 4115 8448 4149 8450
rect 4373 8552 4407 8554
rect 4373 8520 4407 8552
rect 4373 8450 4407 8482
rect 4373 8448 4407 8450
rect 4631 8552 4665 8554
rect 4631 8520 4665 8552
rect 4631 8450 4665 8482
rect 4631 8448 4665 8450
rect 4889 8552 4923 8554
rect 4889 8520 4923 8552
rect 4889 8450 4923 8482
rect 4889 8448 4923 8450
rect 5147 8552 5181 8554
rect 5147 8520 5181 8552
rect 5147 8450 5181 8482
rect 5147 8448 5181 8450
rect 2969 8357 3003 8363
rect 2969 8329 3003 8357
rect 3176 8329 3178 8363
rect 3178 8329 3210 8363
rect 3248 8329 3280 8363
rect 3280 8329 3282 8363
rect 3434 8329 3436 8363
rect 3436 8329 3468 8363
rect 3506 8329 3538 8363
rect 3538 8329 3540 8363
rect 3692 8329 3694 8363
rect 3694 8329 3726 8363
rect 3764 8329 3796 8363
rect 3796 8329 3798 8363
rect 4466 8329 4468 8363
rect 4468 8329 4500 8363
rect 4538 8329 4570 8363
rect 4570 8329 4572 8363
rect 4724 8329 4726 8363
rect 4726 8329 4758 8363
rect 4796 8329 4828 8363
rect 4828 8329 4830 8363
rect 4982 8329 4984 8363
rect 4984 8329 5016 8363
rect 5054 8329 5086 8363
rect 5086 8329 5088 8363
rect 7102 10845 7104 10879
rect 7104 10845 7136 10879
rect 7174 10845 7206 10879
rect 7206 10845 7208 10879
rect 8392 10845 8394 10879
rect 8394 10845 8426 10879
rect 8464 10845 8496 10879
rect 8496 10845 8498 10879
rect 7009 10749 7043 10751
rect 7009 10717 7043 10749
rect 7009 10647 7043 10679
rect 7009 10645 7043 10647
rect 7267 10749 7301 10751
rect 7267 10717 7301 10749
rect 7267 10647 7301 10679
rect 7267 10645 7301 10647
rect 7525 10749 7559 10751
rect 7525 10717 7559 10749
rect 7525 10647 7559 10679
rect 7525 10645 7559 10647
rect 7783 10749 7817 10751
rect 7783 10717 7817 10749
rect 7783 10647 7817 10679
rect 7783 10645 7817 10647
rect 8041 10749 8075 10751
rect 8041 10717 8075 10749
rect 8041 10647 8075 10679
rect 8041 10645 8075 10647
rect 8299 10749 8333 10751
rect 8299 10717 8333 10749
rect 8299 10647 8333 10679
rect 8299 10645 8333 10647
rect 8557 10749 8591 10751
rect 8557 10717 8591 10749
rect 8557 10647 8591 10679
rect 8557 10645 8591 10647
rect 7102 10517 7104 10551
rect 7104 10517 7136 10551
rect 7174 10517 7206 10551
rect 7206 10517 7208 10551
rect 7360 10517 7362 10551
rect 7362 10517 7394 10551
rect 7432 10517 7464 10551
rect 7464 10517 7466 10551
rect 7618 10517 7620 10551
rect 7620 10517 7652 10551
rect 7690 10517 7722 10551
rect 7722 10517 7724 10551
rect 7876 10517 7878 10551
rect 7878 10517 7910 10551
rect 7948 10517 7980 10551
rect 7980 10517 7982 10551
rect 8134 10517 8136 10551
rect 8136 10517 8168 10551
rect 8206 10517 8238 10551
rect 8238 10517 8240 10551
rect 8392 10517 8394 10551
rect 8394 10517 8426 10551
rect 8464 10517 8496 10551
rect 8496 10517 8498 10551
rect 7102 10409 7104 10443
rect 7104 10409 7136 10443
rect 7174 10409 7206 10443
rect 7206 10409 7208 10443
rect 7360 10409 7362 10443
rect 7362 10409 7394 10443
rect 7432 10409 7464 10443
rect 7464 10409 7466 10443
rect 7618 10409 7620 10443
rect 7620 10409 7652 10443
rect 7690 10409 7722 10443
rect 7722 10409 7724 10443
rect 7876 10409 7878 10443
rect 7878 10409 7910 10443
rect 7948 10409 7980 10443
rect 7980 10409 7982 10443
rect 8134 10409 8136 10443
rect 8136 10409 8168 10443
rect 8206 10409 8238 10443
rect 8238 10409 8240 10443
rect 8392 10409 8394 10443
rect 8394 10409 8426 10443
rect 8464 10409 8496 10443
rect 8496 10409 8498 10443
rect 7009 10313 7043 10315
rect 7009 10281 7043 10313
rect 7009 10211 7043 10243
rect 7009 10209 7043 10211
rect 7267 10313 7301 10315
rect 7267 10281 7301 10313
rect 7267 10211 7301 10243
rect 7267 10209 7301 10211
rect 7525 10313 7559 10315
rect 7525 10281 7559 10313
rect 7525 10211 7559 10243
rect 7525 10209 7559 10211
rect 7783 10313 7817 10315
rect 7783 10281 7817 10313
rect 7783 10211 7817 10243
rect 7783 10209 7817 10211
rect 8041 10313 8075 10315
rect 8041 10281 8075 10313
rect 8041 10211 8075 10243
rect 8041 10209 8075 10211
rect 8299 10313 8333 10315
rect 8299 10281 8333 10313
rect 8299 10211 8333 10243
rect 8299 10209 8333 10211
rect 8557 10313 8591 10315
rect 8557 10281 8591 10313
rect 8557 10211 8591 10243
rect 8557 10209 8591 10211
rect 7102 10081 7104 10115
rect 7104 10081 7136 10115
rect 7174 10081 7206 10115
rect 7206 10081 7208 10115
rect 8392 10081 8394 10115
rect 8394 10081 8426 10115
rect 8464 10081 8496 10115
rect 8496 10081 8498 10115
rect 7102 9973 7104 10007
rect 7104 9973 7136 10007
rect 7174 9973 7206 10007
rect 7206 9973 7208 10007
rect 8392 9973 8394 10007
rect 8394 9973 8426 10007
rect 8464 9973 8496 10007
rect 8496 9973 8498 10007
rect 7009 9877 7043 9879
rect 7009 9845 7043 9877
rect 7009 9775 7043 9807
rect 7009 9773 7043 9775
rect 7267 9877 7301 9879
rect 7267 9845 7301 9877
rect 7267 9775 7301 9807
rect 7267 9773 7301 9775
rect 7525 9877 7559 9879
rect 7525 9845 7559 9877
rect 7525 9775 7559 9807
rect 7525 9773 7559 9775
rect 7783 9877 7817 9879
rect 7783 9845 7817 9877
rect 7783 9775 7817 9807
rect 7783 9773 7817 9775
rect 8041 9877 8075 9879
rect 8041 9845 8075 9877
rect 8041 9775 8075 9807
rect 8041 9773 8075 9775
rect 8299 9877 8333 9879
rect 8299 9845 8333 9877
rect 8299 9775 8333 9807
rect 8299 9773 8333 9775
rect 8557 9877 8591 9879
rect 8557 9845 8591 9877
rect 8557 9775 8591 9807
rect 8557 9773 8591 9775
rect 7102 9645 7104 9679
rect 7104 9645 7136 9679
rect 7174 9645 7206 9679
rect 7206 9645 7208 9679
rect 7360 9645 7362 9679
rect 7362 9645 7394 9679
rect 7432 9645 7464 9679
rect 7464 9645 7466 9679
rect 7618 9645 7620 9679
rect 7620 9645 7652 9679
rect 7690 9645 7722 9679
rect 7722 9645 7724 9679
rect 7876 9645 7878 9679
rect 7878 9645 7910 9679
rect 7948 9645 7980 9679
rect 7980 9645 7982 9679
rect 8134 9645 8136 9679
rect 8136 9645 8168 9679
rect 8206 9645 8238 9679
rect 8238 9645 8240 9679
rect 8392 9645 8394 9679
rect 8394 9645 8426 9679
rect 8464 9645 8496 9679
rect 8496 9645 8498 9679
rect 7102 9537 7104 9571
rect 7104 9537 7136 9571
rect 7174 9537 7206 9571
rect 7206 9537 7208 9571
rect 7360 9537 7362 9571
rect 7362 9537 7394 9571
rect 7432 9537 7464 9571
rect 7464 9537 7466 9571
rect 7618 9537 7620 9571
rect 7620 9537 7652 9571
rect 7690 9537 7722 9571
rect 7722 9537 7724 9571
rect 7876 9537 7878 9571
rect 7878 9537 7910 9571
rect 7948 9537 7980 9571
rect 7980 9537 7982 9571
rect 8134 9537 8136 9571
rect 8136 9537 8168 9571
rect 8206 9537 8238 9571
rect 8238 9537 8240 9571
rect 8392 9537 8394 9571
rect 8394 9537 8426 9571
rect 8464 9537 8496 9571
rect 8496 9537 8498 9571
rect 7009 9441 7043 9443
rect 7009 9409 7043 9441
rect 7009 9339 7043 9371
rect 7009 9337 7043 9339
rect 7267 9441 7301 9443
rect 7267 9409 7301 9441
rect 7267 9339 7301 9371
rect 7267 9337 7301 9339
rect 7525 9441 7559 9443
rect 7525 9409 7559 9441
rect 7525 9339 7559 9371
rect 7525 9337 7559 9339
rect 7783 9441 7817 9443
rect 7783 9409 7817 9441
rect 7783 9339 7817 9371
rect 7783 9337 7817 9339
rect 8041 9441 8075 9443
rect 8041 9409 8075 9441
rect 8041 9339 8075 9371
rect 8041 9337 8075 9339
rect 8299 9441 8333 9443
rect 8299 9409 8333 9441
rect 8299 9339 8333 9371
rect 8299 9337 8333 9339
rect 8557 9441 8591 9443
rect 8557 9409 8591 9441
rect 8557 9339 8591 9371
rect 8557 9337 8591 9339
rect 7102 9209 7104 9243
rect 7104 9209 7136 9243
rect 7174 9209 7206 9243
rect 7206 9209 7208 9243
rect 8392 9209 8394 9243
rect 8394 9209 8426 9243
rect 8464 9209 8496 9243
rect 8496 9209 8498 9243
rect 7102 9101 7104 9135
rect 7104 9101 7136 9135
rect 7174 9101 7206 9135
rect 7206 9101 7208 9135
rect 8392 9101 8394 9135
rect 8394 9101 8426 9135
rect 8464 9101 8496 9135
rect 8496 9101 8498 9135
rect 7009 9005 7043 9007
rect 7009 8973 7043 9005
rect 7009 8903 7043 8935
rect 7009 8901 7043 8903
rect 7267 9005 7301 9007
rect 7267 8973 7301 9005
rect 7267 8903 7301 8935
rect 7267 8901 7301 8903
rect 7525 9005 7559 9007
rect 7525 8973 7559 9005
rect 7525 8903 7559 8935
rect 7525 8901 7559 8903
rect 7783 9005 7817 9007
rect 7783 8973 7817 9005
rect 7783 8903 7817 8935
rect 7783 8901 7817 8903
rect 8041 9005 8075 9007
rect 8041 8973 8075 9005
rect 8041 8903 8075 8935
rect 8041 8901 8075 8903
rect 8299 9005 8333 9007
rect 8299 8973 8333 9005
rect 8299 8903 8333 8935
rect 8299 8901 8333 8903
rect 8557 9005 8591 9007
rect 8557 8973 8591 9005
rect 8557 8903 8591 8935
rect 8557 8901 8591 8903
rect 7102 8773 7104 8807
rect 7104 8773 7136 8807
rect 7174 8773 7206 8807
rect 7206 8773 7208 8807
rect 7360 8773 7362 8807
rect 7362 8773 7394 8807
rect 7432 8773 7464 8807
rect 7464 8773 7466 8807
rect 7618 8773 7620 8807
rect 7620 8773 7652 8807
rect 7690 8773 7722 8807
rect 7722 8773 7724 8807
rect 7876 8773 7878 8807
rect 7878 8773 7910 8807
rect 7948 8773 7980 8807
rect 7980 8773 7982 8807
rect 8134 8773 8136 8807
rect 8136 8773 8168 8807
rect 8206 8773 8238 8807
rect 8238 8773 8240 8807
rect 8392 8773 8394 8807
rect 8394 8773 8426 8807
rect 8464 8773 8496 8807
rect 8496 8773 8498 8807
rect 7102 8665 7104 8699
rect 7104 8665 7136 8699
rect 7174 8665 7206 8699
rect 7206 8665 7208 8699
rect 7360 8665 7362 8699
rect 7362 8665 7394 8699
rect 7432 8665 7464 8699
rect 7464 8665 7466 8699
rect 7618 8665 7620 8699
rect 7620 8665 7652 8699
rect 7690 8665 7722 8699
rect 7722 8665 7724 8699
rect 7876 8665 7878 8699
rect 7878 8665 7910 8699
rect 7948 8665 7980 8699
rect 7980 8665 7982 8699
rect 8134 8665 8136 8699
rect 8136 8665 8168 8699
rect 8206 8665 8238 8699
rect 8238 8665 8240 8699
rect 8392 8665 8394 8699
rect 8394 8665 8426 8699
rect 8464 8665 8496 8699
rect 8496 8665 8498 8699
rect 7009 8569 7043 8571
rect 7009 8537 7043 8569
rect 7009 8467 7043 8499
rect 7009 8465 7043 8467
rect 7267 8569 7301 8571
rect 7267 8537 7301 8569
rect 7267 8467 7301 8499
rect 7267 8465 7301 8467
rect 7525 8569 7559 8571
rect 7525 8537 7559 8569
rect 7525 8467 7559 8499
rect 7525 8465 7559 8467
rect 7783 8569 7817 8571
rect 7783 8537 7817 8569
rect 7783 8467 7817 8499
rect 7783 8465 7817 8467
rect 8041 8569 8075 8571
rect 8041 8537 8075 8569
rect 8041 8467 8075 8499
rect 8041 8465 8075 8467
rect 8299 8569 8333 8571
rect 8299 8537 8333 8569
rect 8299 8467 8333 8499
rect 8299 8465 8333 8467
rect 8557 8569 8591 8571
rect 8557 8537 8591 8569
rect 8557 8467 8591 8499
rect 8557 8465 8591 8467
rect 7102 8337 7104 8371
rect 7104 8337 7136 8371
rect 7174 8337 7206 8371
rect 7206 8337 7208 8371
rect 8392 8337 8394 8371
rect 8394 8337 8426 8371
rect 8464 8337 8496 8371
rect 8496 8337 8498 8371
rect 7102 8229 7104 8263
rect 7104 8229 7136 8263
rect 7174 8229 7206 8263
rect 7206 8229 7208 8263
rect 7360 8229 7362 8263
rect 7362 8229 7394 8263
rect 7432 8229 7464 8263
rect 7464 8229 7466 8263
rect 7618 8229 7620 8263
rect 7620 8229 7652 8263
rect 7690 8229 7722 8263
rect 7722 8229 7724 8263
rect 7876 8229 7878 8263
rect 7878 8229 7910 8263
rect 7948 8229 7980 8263
rect 7980 8229 7982 8263
rect 8134 8229 8136 8263
rect 8136 8229 8168 8263
rect 8206 8229 8238 8263
rect 8238 8229 8240 8263
rect 8392 8229 8394 8263
rect 8394 8229 8426 8263
rect 8464 8229 8496 8263
rect 8496 8229 8498 8263
rect -2115 7988 -2113 8022
rect -2113 7988 -2081 8022
rect -2043 7988 -2011 8022
rect -2011 7988 -2009 8022
rect -1857 7988 -1855 8022
rect -1855 7988 -1823 8022
rect -1785 7988 -1753 8022
rect -1753 7988 -1751 8022
rect -1599 7988 -1597 8022
rect -1597 7988 -1565 8022
rect -1527 7988 -1495 8022
rect -1495 7988 -1493 8022
rect -1341 7988 -1339 8022
rect -1339 7988 -1307 8022
rect -1269 7988 -1237 8022
rect -1237 7988 -1235 8022
rect -1083 7988 -1081 8022
rect -1081 7988 -1049 8022
rect -1011 7988 -979 8022
rect -979 7988 -977 8022
rect -825 7988 -823 8022
rect -823 7988 -791 8022
rect -753 7988 -721 8022
rect -721 7988 -719 8022
rect -567 7988 -565 8022
rect -565 7988 -533 8022
rect -495 7988 -463 8022
rect -463 7988 -461 8022
rect -309 7988 -307 8022
rect -307 7988 -275 8022
rect -237 7988 -205 8022
rect -205 7988 -203 8022
rect -51 7988 -49 8022
rect -49 7988 -17 8022
rect 21 7988 53 8022
rect 53 7988 55 8022
rect 207 7988 209 8022
rect 209 7988 241 8022
rect 279 7988 311 8022
rect 311 7988 313 8022
rect 465 7988 467 8022
rect 467 7988 499 8022
rect 537 7988 569 8022
rect 569 7988 571 8022
rect 723 7988 725 8022
rect 725 7988 757 8022
rect 795 7988 827 8022
rect 827 7988 829 8022
rect 981 7988 983 8022
rect 983 7988 1015 8022
rect 1053 7988 1085 8022
rect 1085 7988 1087 8022
rect 1239 7988 1241 8022
rect 1241 7988 1273 8022
rect 1311 7988 1343 8022
rect 1343 7988 1345 8022
rect -2208 7901 -2174 7903
rect -2208 7869 -2174 7901
rect -2208 7799 -2174 7831
rect -2208 7797 -2174 7799
rect -1950 7901 -1916 7903
rect -1950 7869 -1916 7901
rect -1950 7799 -1916 7831
rect -1950 7797 -1916 7799
rect -1692 7901 -1658 7903
rect -1692 7869 -1658 7901
rect -1692 7799 -1658 7831
rect -1692 7797 -1658 7799
rect -1434 7901 -1400 7903
rect -1434 7869 -1400 7901
rect -1434 7799 -1400 7831
rect -1434 7797 -1400 7799
rect -1176 7901 -1142 7903
rect -1176 7869 -1142 7901
rect -1176 7799 -1142 7831
rect -1176 7797 -1142 7799
rect -918 7901 -884 7903
rect -918 7869 -884 7901
rect -918 7799 -884 7831
rect -918 7797 -884 7799
rect -660 7901 -626 7903
rect -660 7869 -626 7901
rect -660 7799 -626 7831
rect -660 7797 -626 7799
rect -402 7901 -368 7903
rect -402 7869 -368 7901
rect -402 7799 -368 7831
rect -402 7797 -368 7799
rect -144 7901 -110 7903
rect -144 7869 -110 7901
rect -144 7799 -110 7831
rect -144 7797 -110 7799
rect 114 7901 148 7903
rect 114 7869 148 7901
rect 114 7799 148 7831
rect 114 7797 148 7799
rect 372 7901 406 7903
rect 372 7869 406 7901
rect 372 7799 406 7831
rect 372 7797 406 7799
rect 630 7901 664 7903
rect 630 7869 664 7901
rect 630 7799 664 7831
rect 630 7797 664 7799
rect 888 7901 922 7903
rect 888 7869 922 7901
rect 888 7799 922 7831
rect 888 7797 922 7799
rect 1146 7901 1180 7903
rect 1146 7869 1180 7901
rect 1146 7799 1180 7831
rect 1146 7797 1180 7799
rect 1404 7901 1438 7903
rect 1404 7869 1438 7901
rect 1404 7799 1438 7831
rect 1404 7797 1438 7799
rect 7009 8133 7043 8135
rect 7009 8101 7043 8133
rect 7009 8031 7043 8063
rect 7009 8029 7043 8031
rect 7267 8133 7301 8135
rect 7267 8101 7301 8133
rect 7267 8031 7301 8063
rect 7267 8029 7301 8031
rect 7525 8133 7559 8135
rect 7525 8101 7559 8133
rect 7525 8031 7559 8063
rect 7525 8029 7559 8031
rect 7783 8133 7817 8135
rect 7783 8101 7817 8133
rect 7783 8031 7817 8063
rect 7783 8029 7817 8031
rect 8041 8133 8075 8135
rect 8041 8101 8075 8133
rect 8041 8031 8075 8063
rect 8041 8029 8075 8031
rect 8299 8133 8333 8135
rect 8299 8101 8333 8133
rect 8299 8031 8333 8063
rect 8299 8029 8333 8031
rect 8557 8133 8591 8135
rect 8557 8101 8591 8133
rect 8557 8031 8591 8063
rect 8557 8029 8591 8031
rect 7102 7901 7104 7935
rect 7104 7901 7136 7935
rect 7174 7901 7206 7935
rect 7206 7901 7208 7935
rect 8392 7901 8394 7935
rect 8394 7901 8426 7935
rect 8464 7901 8496 7935
rect 8496 7901 8498 7935
rect -2115 7678 -2113 7712
rect -2113 7678 -2081 7712
rect -2043 7678 -2011 7712
rect -2011 7678 -2009 7712
rect 1239 7678 1241 7712
rect 1241 7678 1273 7712
rect 1311 7678 1343 7712
rect 1343 7678 1345 7712
rect -2115 7570 -2113 7604
rect -2113 7570 -2081 7604
rect -2043 7570 -2011 7604
rect -2011 7570 -2009 7604
rect -1857 7570 -1855 7604
rect -1855 7570 -1823 7604
rect -1785 7570 -1753 7604
rect -1753 7570 -1751 7604
rect -1599 7570 -1597 7604
rect -1597 7570 -1565 7604
rect -1527 7570 -1495 7604
rect -1495 7570 -1493 7604
rect -1341 7570 -1339 7604
rect -1339 7570 -1307 7604
rect -1269 7570 -1237 7604
rect -1237 7570 -1235 7604
rect -1083 7570 -1081 7604
rect -1081 7570 -1049 7604
rect -1011 7570 -979 7604
rect -979 7570 -977 7604
rect -309 7570 -307 7604
rect -307 7570 -275 7604
rect -237 7570 -205 7604
rect -205 7570 -203 7604
rect -51 7570 -49 7604
rect -49 7570 -17 7604
rect 21 7570 53 7604
rect 53 7570 55 7604
rect 723 7570 725 7604
rect 725 7570 757 7604
rect 795 7570 827 7604
rect 827 7570 829 7604
rect 981 7570 983 7604
rect 983 7570 1015 7604
rect 1053 7570 1085 7604
rect 1085 7570 1087 7604
rect 1239 7570 1241 7604
rect 1241 7570 1273 7604
rect 1311 7570 1343 7604
rect 1343 7570 1345 7604
rect -2208 7483 -2174 7485
rect -2208 7451 -2174 7483
rect -2208 7381 -2174 7413
rect -2208 7379 -2174 7381
rect -1950 7483 -1916 7485
rect -1950 7451 -1916 7483
rect -1950 7381 -1916 7413
rect -1950 7379 -1916 7381
rect -1692 7483 -1658 7485
rect -1692 7451 -1658 7483
rect -1692 7381 -1658 7413
rect -1692 7379 -1658 7381
rect -1434 7483 -1400 7485
rect -1434 7451 -1400 7483
rect -1434 7381 -1400 7413
rect -1434 7379 -1400 7381
rect -1176 7483 -1142 7485
rect -1176 7451 -1142 7483
rect -1176 7381 -1142 7413
rect -1176 7379 -1142 7381
rect -918 7483 -884 7485
rect -918 7451 -884 7483
rect -918 7381 -884 7413
rect -918 7379 -884 7381
rect -660 7483 -626 7485
rect -660 7451 -626 7483
rect -660 7381 -626 7413
rect -660 7379 -626 7381
rect -402 7483 -368 7485
rect -402 7451 -368 7483
rect -402 7381 -368 7413
rect -402 7379 -368 7381
rect -144 7483 -110 7485
rect -144 7451 -110 7483
rect -144 7381 -110 7413
rect -144 7379 -110 7381
rect 114 7483 148 7485
rect 114 7451 148 7483
rect 114 7381 148 7413
rect 114 7379 148 7381
rect 372 7483 406 7485
rect 372 7451 406 7483
rect 372 7381 406 7413
rect 372 7379 406 7381
rect 630 7483 664 7485
rect 630 7451 664 7483
rect 630 7381 664 7413
rect 630 7379 664 7381
rect 888 7483 922 7485
rect 888 7451 922 7483
rect 888 7381 922 7413
rect 888 7379 922 7381
rect 1146 7483 1180 7485
rect 1146 7451 1180 7483
rect 1146 7381 1180 7413
rect 1146 7379 1180 7381
rect 1404 7483 1438 7485
rect 1404 7451 1438 7483
rect 1404 7381 1438 7413
rect 1404 7379 1438 7381
rect 9940 7603 10262 7605
rect 9940 7501 10262 7603
rect 9940 7499 10262 7501
rect -2115 7260 -2113 7294
rect -2113 7260 -2081 7294
rect -2043 7260 -2011 7294
rect -2011 7260 -2009 7294
rect -825 7260 -823 7294
rect -823 7260 -791 7294
rect -753 7260 -721 7294
rect -721 7260 -719 7294
rect -567 7260 -565 7294
rect -565 7260 -533 7294
rect -495 7260 -463 7294
rect -463 7260 -461 7294
rect 207 7260 209 7294
rect 209 7260 241 7294
rect 279 7260 311 7294
rect 311 7260 313 7294
rect 465 7260 467 7294
rect 467 7260 499 7294
rect 537 7260 569 7294
rect 569 7260 571 7294
rect 1239 7260 1241 7294
rect 1241 7260 1273 7294
rect 1311 7260 1343 7294
rect 1343 7260 1345 7294
rect -2115 7152 -2113 7186
rect -2113 7152 -2081 7186
rect -2043 7152 -2011 7186
rect -2011 7152 -2009 7186
rect -1857 7152 -1855 7186
rect -1855 7152 -1823 7186
rect -1785 7152 -1753 7186
rect -1753 7152 -1751 7186
rect -1599 7152 -1597 7186
rect -1597 7152 -1565 7186
rect -1527 7152 -1495 7186
rect -1495 7152 -1493 7186
rect -825 7152 -823 7186
rect -823 7152 -791 7186
rect -753 7152 -721 7186
rect -721 7152 -719 7186
rect -567 7152 -565 7186
rect -565 7152 -533 7186
rect -495 7152 -463 7186
rect -463 7152 -461 7186
rect 207 7152 209 7186
rect 209 7152 241 7186
rect 279 7152 311 7186
rect 311 7152 313 7186
rect 465 7152 467 7186
rect 467 7152 499 7186
rect 537 7152 569 7186
rect 569 7152 571 7186
rect 1239 7152 1241 7186
rect 1241 7152 1273 7186
rect 1311 7152 1343 7186
rect 1343 7152 1345 7186
rect -2208 7065 -2174 7067
rect -2208 7033 -2174 7065
rect -2208 6963 -2174 6995
rect -2208 6961 -2174 6963
rect -1950 7065 -1916 7067
rect -1950 7033 -1916 7065
rect -1950 6963 -1916 6995
rect -1950 6961 -1916 6963
rect -1692 7065 -1658 7067
rect -1692 7033 -1658 7065
rect -1692 6963 -1658 6995
rect -1692 6961 -1658 6963
rect -1434 7065 -1400 7067
rect -1434 7033 -1400 7065
rect -1434 6963 -1400 6995
rect -1434 6961 -1400 6963
rect -1176 7065 -1142 7067
rect -1176 7033 -1142 7065
rect -1176 6963 -1142 6995
rect -1176 6961 -1142 6963
rect -918 7065 -884 7067
rect -918 7033 -884 7065
rect -918 6963 -884 6995
rect -918 6961 -884 6963
rect -660 7065 -626 7067
rect -660 7033 -626 7065
rect -660 6963 -626 6995
rect -660 6961 -626 6963
rect -402 7065 -368 7067
rect -402 7033 -368 7065
rect -402 6963 -368 6995
rect -402 6961 -368 6963
rect -144 7065 -110 7067
rect -144 7033 -110 7065
rect -144 6963 -110 6995
rect -144 6961 -110 6963
rect 114 7065 148 7067
rect 114 7033 148 7065
rect 114 6963 148 6995
rect 114 6961 148 6963
rect 372 7065 406 7067
rect 372 7033 406 7065
rect 372 6963 406 6995
rect 372 6961 406 6963
rect 630 7065 664 7067
rect 630 7033 664 7065
rect 630 6963 664 6995
rect 630 6961 664 6963
rect 888 7065 922 7067
rect 888 7033 922 7065
rect 888 6963 922 6995
rect 888 6961 922 6963
rect 1146 7065 1180 7067
rect 1146 7033 1180 7065
rect 1146 6963 1180 6995
rect 1146 6961 1180 6963
rect 1404 7065 1438 7067
rect 1404 7033 1438 7065
rect 1404 6963 1438 6995
rect 1404 6961 1438 6963
rect -2115 6842 -2113 6876
rect -2113 6842 -2081 6876
rect -2043 6842 -2011 6876
rect -2011 6842 -2009 6876
rect -1341 6842 -1339 6876
rect -1339 6842 -1307 6876
rect -1269 6842 -1237 6876
rect -1237 6842 -1235 6876
rect -1083 6842 -1081 6876
rect -1081 6842 -1049 6876
rect -1011 6842 -979 6876
rect -979 6842 -977 6876
rect -309 6842 -307 6876
rect -307 6842 -275 6876
rect -237 6842 -205 6876
rect -205 6842 -203 6876
rect -51 6842 -49 6876
rect -49 6842 -17 6876
rect 21 6842 53 6876
rect 53 6842 55 6876
rect 723 6842 725 6876
rect 725 6842 757 6876
rect 795 6842 827 6876
rect 827 6842 829 6876
rect 981 6842 983 6876
rect 983 6842 1015 6876
rect 1053 6842 1085 6876
rect 1085 6842 1087 6876
rect 1239 6842 1241 6876
rect 1241 6842 1273 6876
rect 1311 6842 1343 6876
rect 1343 6842 1345 6876
rect -2115 6734 -2113 6768
rect -2113 6734 -2081 6768
rect -2043 6734 -2011 6768
rect -2011 6734 -2009 6768
rect -1341 6734 -1339 6768
rect -1339 6734 -1307 6768
rect -1269 6734 -1237 6768
rect -1237 6734 -1235 6768
rect -1083 6734 -1081 6768
rect -1081 6734 -1049 6768
rect -1011 6734 -979 6768
rect -979 6734 -977 6768
rect -309 6734 -307 6768
rect -307 6734 -275 6768
rect -237 6734 -205 6768
rect -205 6734 -203 6768
rect -51 6734 -49 6768
rect -49 6734 -17 6768
rect 21 6734 53 6768
rect 53 6734 55 6768
rect 723 6734 725 6768
rect 725 6734 757 6768
rect 795 6734 827 6768
rect 827 6734 829 6768
rect 981 6734 983 6768
rect 983 6734 1015 6768
rect 1053 6734 1085 6768
rect 1085 6734 1087 6768
rect 1239 6734 1241 6768
rect 1241 6734 1273 6768
rect 1311 6734 1343 6768
rect 1343 6734 1345 6768
rect -2208 6647 -2174 6649
rect -2208 6615 -2174 6647
rect -2208 6545 -2174 6577
rect -2208 6543 -2174 6545
rect -1950 6647 -1916 6649
rect -1950 6615 -1916 6647
rect -1950 6545 -1916 6577
rect -1950 6543 -1916 6545
rect -1692 6647 -1658 6649
rect -1692 6615 -1658 6647
rect -1692 6545 -1658 6577
rect -1692 6543 -1658 6545
rect -1434 6647 -1400 6649
rect -1434 6615 -1400 6647
rect -1434 6545 -1400 6577
rect -1434 6543 -1400 6545
rect -1176 6647 -1142 6649
rect -1176 6615 -1142 6647
rect -1176 6545 -1142 6577
rect -1176 6543 -1142 6545
rect -918 6647 -884 6649
rect -918 6615 -884 6647
rect -918 6545 -884 6577
rect -918 6543 -884 6545
rect -660 6647 -626 6649
rect -660 6615 -626 6647
rect -660 6545 -626 6577
rect -660 6543 -626 6545
rect -402 6647 -368 6649
rect -402 6615 -368 6647
rect -402 6545 -368 6577
rect -402 6543 -368 6545
rect -144 6647 -110 6649
rect -144 6615 -110 6647
rect -144 6545 -110 6577
rect -144 6543 -110 6545
rect 114 6647 148 6649
rect 114 6615 148 6647
rect 114 6545 148 6577
rect 114 6543 148 6545
rect 372 6647 406 6649
rect 372 6615 406 6647
rect 372 6545 406 6577
rect 372 6543 406 6545
rect 630 6647 664 6649
rect 630 6615 664 6647
rect 630 6545 664 6577
rect 630 6543 664 6545
rect 888 6647 922 6649
rect 888 6615 922 6647
rect 888 6545 922 6577
rect 888 6543 922 6545
rect 1146 6647 1180 6649
rect 1146 6615 1180 6647
rect 1146 6545 1180 6577
rect 1146 6543 1180 6545
rect 1404 6647 1438 6649
rect 1404 6615 1438 6647
rect 1404 6545 1438 6577
rect 1404 6543 1438 6545
rect -2115 6424 -2113 6458
rect -2113 6424 -2081 6458
rect -2043 6424 -2011 6458
rect -2011 6424 -2009 6458
rect -1857 6424 -1855 6458
rect -1855 6424 -1823 6458
rect -1785 6424 -1753 6458
rect -1753 6424 -1751 6458
rect -1599 6424 -1597 6458
rect -1597 6424 -1565 6458
rect -1527 6424 -1495 6458
rect -1495 6424 -1493 6458
rect -825 6424 -823 6458
rect -823 6424 -791 6458
rect -753 6424 -721 6458
rect -721 6424 -719 6458
rect -567 6424 -565 6458
rect -565 6424 -533 6458
rect -495 6424 -463 6458
rect -463 6424 -461 6458
rect 207 6424 209 6458
rect 209 6424 241 6458
rect 279 6424 311 6458
rect 311 6424 313 6458
rect 465 6424 467 6458
rect 467 6424 499 6458
rect 537 6424 569 6458
rect 569 6424 571 6458
rect 1239 6424 1241 6458
rect 1241 6424 1273 6458
rect 1311 6424 1343 6458
rect 1343 6424 1345 6458
rect -2115 6316 -2113 6350
rect -2113 6316 -2081 6350
rect -2043 6316 -2011 6350
rect -2011 6316 -2009 6350
rect -1857 6316 -1855 6350
rect -1855 6316 -1823 6350
rect -1785 6316 -1753 6350
rect -1753 6316 -1751 6350
rect -1599 6316 -1597 6350
rect -1597 6316 -1565 6350
rect -1527 6316 -1495 6350
rect -1495 6316 -1493 6350
rect -825 6316 -823 6350
rect -823 6316 -791 6350
rect -753 6316 -721 6350
rect -721 6316 -719 6350
rect -567 6316 -565 6350
rect -565 6316 -533 6350
rect -495 6316 -463 6350
rect -463 6316 -461 6350
rect 207 6316 209 6350
rect 209 6316 241 6350
rect 279 6316 311 6350
rect 311 6316 313 6350
rect 465 6316 467 6350
rect 467 6316 499 6350
rect 537 6316 569 6350
rect 569 6316 571 6350
rect 1239 6316 1241 6350
rect 1241 6316 1273 6350
rect 1311 6316 1343 6350
rect 1343 6316 1345 6350
rect -2208 6229 -2174 6231
rect -2208 6197 -2174 6229
rect -2208 6127 -2174 6159
rect -2208 6125 -2174 6127
rect -1950 6229 -1916 6231
rect -1950 6197 -1916 6229
rect -1950 6127 -1916 6159
rect -1950 6125 -1916 6127
rect -1692 6229 -1658 6231
rect -1692 6197 -1658 6229
rect -1692 6127 -1658 6159
rect -1692 6125 -1658 6127
rect -1434 6229 -1400 6231
rect -1434 6197 -1400 6229
rect -1434 6127 -1400 6159
rect -1434 6125 -1400 6127
rect -1176 6229 -1142 6231
rect -1176 6197 -1142 6229
rect -1176 6127 -1142 6159
rect -1176 6125 -1142 6127
rect -918 6229 -884 6231
rect -918 6197 -884 6229
rect -918 6127 -884 6159
rect -918 6125 -884 6127
rect -660 6229 -626 6231
rect -660 6197 -626 6229
rect -660 6127 -626 6159
rect -660 6125 -626 6127
rect -402 6229 -368 6231
rect -402 6197 -368 6229
rect -402 6127 -368 6159
rect -402 6125 -368 6127
rect -144 6229 -110 6231
rect -144 6197 -110 6229
rect -144 6127 -110 6159
rect -144 6125 -110 6127
rect 114 6229 148 6231
rect 114 6197 148 6229
rect 114 6127 148 6159
rect 114 6125 148 6127
rect 372 6229 406 6231
rect 372 6197 406 6229
rect 372 6127 406 6159
rect 372 6125 406 6127
rect 630 6229 664 6231
rect 630 6197 664 6229
rect 630 6127 664 6159
rect 630 6125 664 6127
rect 888 6229 922 6231
rect 888 6197 922 6229
rect 888 6127 922 6159
rect 888 6125 922 6127
rect 1146 6229 1180 6231
rect 1146 6197 1180 6229
rect 1146 6127 1180 6159
rect 1146 6125 1180 6127
rect 1404 6229 1438 6231
rect 1404 6197 1438 6229
rect 1404 6127 1438 6159
rect 1404 6125 1438 6127
rect -2115 6006 -2113 6040
rect -2113 6006 -2081 6040
rect -2043 6006 -2011 6040
rect -2011 6006 -2009 6040
rect -1341 6006 -1339 6040
rect -1339 6006 -1307 6040
rect -1269 6006 -1237 6040
rect -1237 6006 -1235 6040
rect -1083 6006 -1081 6040
rect -1081 6006 -1049 6040
rect -1011 6006 -979 6040
rect -979 6006 -977 6040
rect -309 6006 -307 6040
rect -307 6006 -275 6040
rect -237 6006 -205 6040
rect -205 6006 -203 6040
rect -51 6006 -49 6040
rect -49 6006 -17 6040
rect 21 6006 53 6040
rect 53 6006 55 6040
rect 723 6006 725 6040
rect 725 6006 757 6040
rect 795 6006 827 6040
rect 827 6006 829 6040
rect 981 6006 983 6040
rect 983 6006 1015 6040
rect 1053 6006 1085 6040
rect 1085 6006 1087 6040
rect 1239 6006 1241 6040
rect 1241 6006 1273 6040
rect 1311 6006 1343 6040
rect 1343 6006 1345 6040
rect -2115 5898 -2113 5932
rect -2113 5898 -2081 5932
rect -2043 5898 -2011 5932
rect -2011 5898 -2009 5932
rect -1341 5898 -1339 5932
rect -1339 5898 -1307 5932
rect -1269 5898 -1237 5932
rect -1237 5898 -1235 5932
rect -1083 5898 -1081 5932
rect -1081 5898 -1049 5932
rect -1011 5898 -979 5932
rect -979 5898 -977 5932
rect -309 5898 -307 5932
rect -307 5898 -275 5932
rect -237 5898 -205 5932
rect -205 5898 -203 5932
rect -51 5898 -49 5932
rect -49 5898 -17 5932
rect 21 5898 53 5932
rect 53 5898 55 5932
rect 723 5898 725 5932
rect 725 5898 757 5932
rect 795 5898 827 5932
rect 827 5898 829 5932
rect 981 5898 983 5932
rect 983 5898 1015 5932
rect 1053 5898 1085 5932
rect 1085 5898 1087 5932
rect 1239 5898 1241 5932
rect 1241 5898 1273 5932
rect 1311 5898 1343 5932
rect 1343 5898 1345 5932
rect -2208 5811 -2174 5813
rect -2208 5779 -2174 5811
rect -2208 5709 -2174 5741
rect -2208 5707 -2174 5709
rect -1950 5811 -1916 5813
rect -1950 5779 -1916 5811
rect -1950 5709 -1916 5741
rect -1950 5707 -1916 5709
rect -1692 5811 -1658 5813
rect -1692 5779 -1658 5811
rect -1692 5709 -1658 5741
rect -1692 5707 -1658 5709
rect -1434 5811 -1400 5813
rect -1434 5779 -1400 5811
rect -1434 5709 -1400 5741
rect -1434 5707 -1400 5709
rect -1176 5811 -1142 5813
rect -1176 5779 -1142 5811
rect -1176 5709 -1142 5741
rect -1176 5707 -1142 5709
rect -918 5811 -884 5813
rect -918 5779 -884 5811
rect -918 5709 -884 5741
rect -918 5707 -884 5709
rect -660 5811 -626 5813
rect -660 5779 -626 5811
rect -660 5709 -626 5741
rect -660 5707 -626 5709
rect -402 5811 -368 5813
rect -402 5779 -368 5811
rect -402 5709 -368 5741
rect -402 5707 -368 5709
rect -144 5811 -110 5813
rect -144 5779 -110 5811
rect -144 5709 -110 5741
rect -144 5707 -110 5709
rect 114 5811 148 5813
rect 114 5779 148 5811
rect 114 5709 148 5741
rect 114 5707 148 5709
rect 372 5811 406 5813
rect 372 5779 406 5811
rect 372 5709 406 5741
rect 372 5707 406 5709
rect 630 5811 664 5813
rect 630 5779 664 5811
rect 630 5709 664 5741
rect 630 5707 664 5709
rect 888 5811 922 5813
rect 888 5779 922 5811
rect 888 5709 922 5741
rect 888 5707 922 5709
rect 1146 5811 1180 5813
rect 1146 5779 1180 5811
rect 1146 5709 1180 5741
rect 1146 5707 1180 5709
rect 1404 5811 1438 5813
rect 1404 5779 1438 5811
rect 1404 5709 1438 5741
rect 1404 5707 1438 5709
rect -2115 5588 -2113 5622
rect -2113 5588 -2081 5622
rect -2043 5588 -2011 5622
rect -2011 5588 -2009 5622
rect -1857 5588 -1855 5622
rect -1855 5588 -1823 5622
rect -1785 5588 -1753 5622
rect -1753 5588 -1751 5622
rect -1599 5588 -1597 5622
rect -1597 5588 -1565 5622
rect -1527 5588 -1495 5622
rect -1495 5588 -1493 5622
rect -825 5588 -823 5622
rect -823 5588 -791 5622
rect -753 5588 -721 5622
rect -721 5588 -719 5622
rect -567 5588 -565 5622
rect -565 5588 -533 5622
rect -495 5588 -463 5622
rect -463 5588 -461 5622
rect 207 5588 209 5622
rect 209 5588 241 5622
rect 279 5588 311 5622
rect 311 5588 313 5622
rect 465 5588 467 5622
rect 467 5588 499 5622
rect 537 5588 569 5622
rect 569 5588 571 5622
rect 1239 5588 1241 5622
rect 1241 5588 1273 5622
rect 1311 5588 1343 5622
rect 1343 5588 1345 5622
rect -2115 5480 -2113 5514
rect -2113 5480 -2081 5514
rect -2043 5480 -2011 5514
rect -2011 5480 -2009 5514
rect -1857 5480 -1855 5514
rect -1855 5480 -1823 5514
rect -1785 5480 -1753 5514
rect -1753 5480 -1751 5514
rect -1599 5480 -1597 5514
rect -1597 5480 -1565 5514
rect -1527 5480 -1495 5514
rect -1495 5480 -1493 5514
rect -825 5480 -823 5514
rect -823 5480 -791 5514
rect -753 5480 -721 5514
rect -721 5480 -719 5514
rect -567 5480 -565 5514
rect -565 5480 -533 5514
rect -495 5480 -463 5514
rect -463 5480 -461 5514
rect 207 5480 209 5514
rect 209 5480 241 5514
rect 279 5480 311 5514
rect 311 5480 313 5514
rect 465 5480 467 5514
rect 467 5480 499 5514
rect 537 5480 569 5514
rect 569 5480 571 5514
rect 1239 5480 1241 5514
rect 1241 5480 1273 5514
rect 1311 5480 1343 5514
rect 1343 5480 1345 5514
rect -2208 5393 -2174 5395
rect -2208 5361 -2174 5393
rect -2208 5291 -2174 5323
rect -2208 5289 -2174 5291
rect -1950 5393 -1916 5395
rect -1950 5361 -1916 5393
rect -1950 5291 -1916 5323
rect -1950 5289 -1916 5291
rect -1692 5393 -1658 5395
rect -1692 5361 -1658 5393
rect -1692 5291 -1658 5323
rect -1692 5289 -1658 5291
rect -1434 5393 -1400 5395
rect -1434 5361 -1400 5393
rect -1434 5291 -1400 5323
rect -1434 5289 -1400 5291
rect -1176 5393 -1142 5395
rect -1176 5361 -1142 5393
rect -1176 5291 -1142 5323
rect -1176 5289 -1142 5291
rect -918 5393 -884 5395
rect -918 5361 -884 5393
rect -918 5291 -884 5323
rect -918 5289 -884 5291
rect -660 5393 -626 5395
rect -660 5361 -626 5393
rect -660 5291 -626 5323
rect -660 5289 -626 5291
rect -402 5393 -368 5395
rect -402 5361 -368 5393
rect -402 5291 -368 5323
rect -402 5289 -368 5291
rect -144 5393 -110 5395
rect -144 5361 -110 5393
rect -144 5291 -110 5323
rect -144 5289 -110 5291
rect 114 5393 148 5395
rect 114 5361 148 5393
rect 114 5291 148 5323
rect 114 5289 148 5291
rect 372 5393 406 5395
rect 372 5361 406 5393
rect 372 5291 406 5323
rect 372 5289 406 5291
rect 630 5393 664 5395
rect 630 5361 664 5393
rect 630 5291 664 5323
rect 630 5289 664 5291
rect 888 5393 922 5395
rect 888 5361 922 5393
rect 888 5291 922 5323
rect 888 5289 922 5291
rect 1146 5393 1180 5395
rect 1146 5361 1180 5393
rect 1146 5291 1180 5323
rect 1146 5289 1180 5291
rect 1404 5393 1438 5395
rect 1404 5361 1438 5393
rect 1404 5291 1438 5323
rect 1404 5289 1438 5291
rect -2115 5170 -2113 5204
rect -2113 5170 -2081 5204
rect -2043 5170 -2011 5204
rect -2011 5170 -2009 5204
rect -1341 5170 -1339 5204
rect -1339 5170 -1307 5204
rect -1269 5170 -1237 5204
rect -1237 5170 -1235 5204
rect -1083 5170 -1081 5204
rect -1081 5170 -1049 5204
rect -1011 5170 -979 5204
rect -979 5170 -977 5204
rect -309 5170 -307 5204
rect -307 5170 -275 5204
rect -237 5170 -205 5204
rect -205 5170 -203 5204
rect -51 5170 -49 5204
rect -49 5170 -17 5204
rect 21 5170 53 5204
rect 53 5170 55 5204
rect 723 5170 725 5204
rect 725 5170 757 5204
rect 795 5170 827 5204
rect 827 5170 829 5204
rect 981 5170 983 5204
rect 983 5170 1015 5204
rect 1053 5170 1085 5204
rect 1085 5170 1087 5204
rect 1239 5170 1241 5204
rect 1241 5170 1273 5204
rect 1311 5170 1343 5204
rect 1343 5170 1345 5204
rect -2115 5062 -2113 5096
rect -2113 5062 -2081 5096
rect -2043 5062 -2011 5096
rect -2011 5062 -2009 5096
rect -1341 5062 -1339 5096
rect -1339 5062 -1307 5096
rect -1269 5062 -1237 5096
rect -1237 5062 -1235 5096
rect -1083 5062 -1081 5096
rect -1081 5062 -1049 5096
rect -1011 5062 -979 5096
rect -979 5062 -977 5096
rect -309 5062 -307 5096
rect -307 5062 -275 5096
rect -237 5062 -205 5096
rect -205 5062 -203 5096
rect -51 5062 -49 5096
rect -49 5062 -17 5096
rect 21 5062 53 5096
rect 53 5062 55 5096
rect 723 5062 725 5096
rect 725 5062 757 5096
rect 795 5062 827 5096
rect 827 5062 829 5096
rect 981 5062 983 5096
rect 983 5062 1015 5096
rect 1053 5062 1085 5096
rect 1085 5062 1087 5096
rect 1239 5062 1241 5096
rect 1241 5062 1273 5096
rect 1311 5062 1343 5096
rect 1343 5062 1345 5096
rect -2208 4975 -2174 4977
rect -2208 4943 -2174 4975
rect -2208 4873 -2174 4905
rect -2208 4871 -2174 4873
rect -1950 4975 -1916 4977
rect -1950 4943 -1916 4975
rect -1950 4873 -1916 4905
rect -1950 4871 -1916 4873
rect -1692 4975 -1658 4977
rect -1692 4943 -1658 4975
rect -1692 4873 -1658 4905
rect -1692 4871 -1658 4873
rect -1434 4975 -1400 4977
rect -1434 4943 -1400 4975
rect -1434 4873 -1400 4905
rect -1434 4871 -1400 4873
rect -1176 4975 -1142 4977
rect -1176 4943 -1142 4975
rect -1176 4873 -1142 4905
rect -1176 4871 -1142 4873
rect -918 4975 -884 4977
rect -918 4943 -884 4975
rect -918 4873 -884 4905
rect -918 4871 -884 4873
rect -660 4975 -626 4977
rect -660 4943 -626 4975
rect -660 4873 -626 4905
rect -660 4871 -626 4873
rect -402 4975 -368 4977
rect -402 4943 -368 4975
rect -402 4873 -368 4905
rect -402 4871 -368 4873
rect -144 4975 -110 4977
rect -144 4943 -110 4975
rect -144 4873 -110 4905
rect -144 4871 -110 4873
rect 114 4975 148 4977
rect 114 4943 148 4975
rect 114 4873 148 4905
rect 114 4871 148 4873
rect 372 4975 406 4977
rect 372 4943 406 4975
rect 372 4873 406 4905
rect 372 4871 406 4873
rect 630 4975 664 4977
rect 630 4943 664 4975
rect 630 4873 664 4905
rect 630 4871 664 4873
rect 888 4975 922 4977
rect 888 4943 922 4975
rect 888 4873 922 4905
rect 888 4871 922 4873
rect 1146 4975 1180 4977
rect 1146 4943 1180 4975
rect 1146 4873 1180 4905
rect 1146 4871 1180 4873
rect 1404 4975 1438 4977
rect 1404 4943 1438 4975
rect 1404 4873 1438 4905
rect 1404 4871 1438 4873
rect -2115 4752 -2113 4786
rect -2113 4752 -2081 4786
rect -2043 4752 -2011 4786
rect -2011 4752 -2009 4786
rect -1857 4752 -1855 4786
rect -1855 4752 -1823 4786
rect -1785 4752 -1753 4786
rect -1753 4752 -1751 4786
rect -1599 4752 -1597 4786
rect -1597 4752 -1565 4786
rect -1527 4752 -1495 4786
rect -1495 4752 -1493 4786
rect -825 4752 -823 4786
rect -823 4752 -791 4786
rect -753 4752 -721 4786
rect -721 4752 -719 4786
rect -567 4752 -565 4786
rect -565 4752 -533 4786
rect -495 4752 -463 4786
rect -463 4752 -461 4786
rect 207 4752 209 4786
rect 209 4752 241 4786
rect 279 4752 311 4786
rect 311 4752 313 4786
rect 465 4752 467 4786
rect 467 4752 499 4786
rect 537 4752 569 4786
rect 569 4752 571 4786
rect 1239 4752 1241 4786
rect 1241 4752 1273 4786
rect 1311 4752 1343 4786
rect 1343 4752 1345 4786
rect -2115 4644 -2113 4678
rect -2113 4644 -2081 4678
rect -2043 4644 -2011 4678
rect -2011 4644 -2009 4678
rect -1857 4644 -1855 4678
rect -1855 4644 -1823 4678
rect -1785 4644 -1753 4678
rect -1753 4644 -1751 4678
rect -1599 4644 -1597 4678
rect -1597 4644 -1565 4678
rect -1527 4644 -1495 4678
rect -1495 4644 -1493 4678
rect -825 4644 -823 4678
rect -823 4644 -791 4678
rect -753 4644 -721 4678
rect -721 4644 -719 4678
rect -567 4644 -565 4678
rect -565 4644 -533 4678
rect -495 4644 -463 4678
rect -463 4644 -461 4678
rect 207 4644 209 4678
rect 209 4644 241 4678
rect 279 4644 311 4678
rect 311 4644 313 4678
rect 465 4644 467 4678
rect 467 4644 499 4678
rect 537 4644 569 4678
rect 569 4644 571 4678
rect 723 4644 725 4678
rect 725 4644 757 4678
rect 795 4644 827 4678
rect 827 4644 829 4678
rect 981 4644 983 4678
rect 983 4644 1015 4678
rect 1053 4644 1085 4678
rect 1085 4644 1087 4678
rect 1239 4644 1241 4678
rect 1241 4644 1273 4678
rect 1311 4644 1343 4678
rect 1343 4644 1345 4678
rect -2208 4557 -2174 4559
rect -2208 4525 -2174 4557
rect -2208 4455 -2174 4487
rect -2208 4453 -2174 4455
rect -1950 4557 -1916 4559
rect -1950 4525 -1916 4557
rect -1950 4455 -1916 4487
rect -1950 4453 -1916 4455
rect -1692 4557 -1658 4559
rect -1692 4525 -1658 4557
rect -1692 4455 -1658 4487
rect -1692 4453 -1658 4455
rect -1434 4557 -1400 4559
rect -1434 4525 -1400 4557
rect -1434 4455 -1400 4487
rect -1434 4453 -1400 4455
rect -1176 4557 -1142 4559
rect -1176 4525 -1142 4557
rect -1176 4455 -1142 4487
rect -1176 4453 -1142 4455
rect -918 4557 -884 4559
rect -918 4525 -884 4557
rect -918 4455 -884 4487
rect -918 4453 -884 4455
rect -660 4557 -626 4559
rect -660 4525 -626 4557
rect -660 4455 -626 4487
rect -660 4453 -626 4455
rect -402 4557 -368 4559
rect -402 4525 -368 4557
rect -402 4455 -368 4487
rect -402 4453 -368 4455
rect -144 4557 -110 4559
rect -144 4525 -110 4557
rect -144 4455 -110 4487
rect -144 4453 -110 4455
rect 114 4557 148 4559
rect 114 4525 148 4557
rect 114 4455 148 4487
rect 114 4453 148 4455
rect 372 4557 406 4559
rect 372 4525 406 4557
rect 372 4455 406 4487
rect 372 4453 406 4455
rect 630 4557 664 4559
rect 630 4525 664 4557
rect 630 4455 664 4487
rect 630 4453 664 4455
rect 888 4557 922 4559
rect 888 4525 922 4557
rect 888 4455 922 4487
rect 888 4453 922 4455
rect 1146 4557 1180 4559
rect 1146 4525 1180 4557
rect 1146 4455 1180 4487
rect 1146 4453 1180 4455
rect 1404 4557 1438 4559
rect 1404 4525 1438 4557
rect 1404 4455 1438 4487
rect 1404 4453 1438 4455
rect -2115 4334 -2113 4368
rect -2113 4334 -2081 4368
rect -2043 4334 -2011 4368
rect -2011 4334 -2009 4368
rect -1341 4334 -1339 4368
rect -1339 4334 -1307 4368
rect -1269 4334 -1237 4368
rect -1237 4334 -1235 4368
rect -1083 4334 -1081 4368
rect -1081 4334 -1049 4368
rect -1011 4334 -979 4368
rect -979 4334 -977 4368
rect -309 4334 -307 4368
rect -307 4334 -275 4368
rect -237 4334 -205 4368
rect -205 4334 -203 4368
rect -51 4334 -49 4368
rect -49 4334 -17 4368
rect 21 4334 53 4368
rect 53 4334 55 4368
rect 1239 4334 1241 4368
rect 1241 4334 1273 4368
rect 1311 4334 1343 4368
rect 1343 4334 1345 4368
rect -2115 4226 -2113 4260
rect -2113 4226 -2081 4260
rect -2043 4226 -2011 4260
rect -2011 4226 -2009 4260
rect -1857 4226 -1855 4260
rect -1855 4226 -1823 4260
rect -1785 4226 -1753 4260
rect -1753 4226 -1751 4260
rect -1599 4226 -1597 4260
rect -1597 4226 -1565 4260
rect -1527 4226 -1495 4260
rect -1495 4226 -1493 4260
rect -1341 4226 -1339 4260
rect -1339 4226 -1307 4260
rect -1269 4226 -1237 4260
rect -1237 4226 -1235 4260
rect -1083 4226 -1081 4260
rect -1081 4226 -1049 4260
rect -1011 4226 -979 4260
rect -979 4226 -977 4260
rect -825 4226 -823 4260
rect -823 4226 -791 4260
rect -753 4226 -721 4260
rect -721 4226 -719 4260
rect -567 4226 -565 4260
rect -565 4226 -533 4260
rect -495 4226 -463 4260
rect -463 4226 -461 4260
rect -309 4226 -307 4260
rect -307 4226 -275 4260
rect -237 4226 -205 4260
rect -205 4226 -203 4260
rect -51 4226 -49 4260
rect -49 4226 -17 4260
rect 21 4226 53 4260
rect 53 4226 55 4260
rect 207 4226 209 4260
rect 209 4226 241 4260
rect 279 4226 311 4260
rect 311 4226 313 4260
rect 465 4226 467 4260
rect 467 4226 499 4260
rect 537 4226 569 4260
rect 569 4226 571 4260
rect 723 4226 725 4260
rect 725 4226 757 4260
rect 795 4226 827 4260
rect 827 4226 829 4260
rect 981 4226 983 4260
rect 983 4226 1015 4260
rect 1053 4226 1085 4260
rect 1085 4226 1087 4260
rect 1239 4226 1241 4260
rect 1241 4226 1273 4260
rect 1311 4226 1343 4260
rect 1343 4226 1345 4260
rect -2208 4139 -2174 4141
rect -2208 4107 -2174 4139
rect -2208 4037 -2174 4069
rect -2208 4035 -2174 4037
rect -1950 4139 -1916 4141
rect -1950 4107 -1916 4139
rect -1950 4037 -1916 4069
rect -1950 4035 -1916 4037
rect -1692 4139 -1658 4141
rect -1692 4107 -1658 4139
rect -1692 4037 -1658 4069
rect -1692 4035 -1658 4037
rect -1434 4139 -1400 4141
rect -1434 4107 -1400 4139
rect -1434 4037 -1400 4069
rect -1434 4035 -1400 4037
rect -1176 4139 -1142 4141
rect -1176 4107 -1142 4139
rect -1176 4037 -1142 4069
rect -1176 4035 -1142 4037
rect -918 4139 -884 4141
rect -918 4107 -884 4139
rect -918 4037 -884 4069
rect -918 4035 -884 4037
rect -660 4139 -626 4141
rect -660 4107 -626 4139
rect -660 4037 -626 4069
rect -660 4035 -626 4037
rect -402 4139 -368 4141
rect -402 4107 -368 4139
rect -402 4037 -368 4069
rect -402 4035 -368 4037
rect -144 4139 -110 4141
rect -144 4107 -110 4139
rect -144 4037 -110 4069
rect -144 4035 -110 4037
rect 114 4139 148 4141
rect 114 4107 148 4139
rect 114 4037 148 4069
rect 114 4035 148 4037
rect 372 4139 406 4141
rect 372 4107 406 4139
rect 372 4037 406 4069
rect 372 4035 406 4037
rect 630 4139 664 4141
rect 630 4107 664 4139
rect 630 4037 664 4069
rect 630 4035 664 4037
rect 888 4139 922 4141
rect 888 4107 922 4139
rect 888 4037 922 4069
rect 888 4035 922 4037
rect 1146 4139 1180 4141
rect 1146 4107 1180 4139
rect 1146 4037 1180 4069
rect 1146 4035 1180 4037
rect 1404 4139 1438 4141
rect 1404 4107 1438 4139
rect 1404 4037 1438 4069
rect 1404 4035 1438 4037
rect 1518 4024 1552 4041
rect 1518 4007 1552 4024
rect 3715 7349 3717 7383
rect 3717 7349 3749 7383
rect 3787 7349 3819 7383
rect 3819 7349 3821 7383
rect 3973 7349 3975 7383
rect 3975 7349 4007 7383
rect 4045 7349 4077 7383
rect 4077 7349 4079 7383
rect 4231 7349 4233 7383
rect 4233 7349 4265 7383
rect 4303 7349 4335 7383
rect 4335 7349 4337 7383
rect 4489 7349 4491 7383
rect 4491 7349 4523 7383
rect 4561 7349 4593 7383
rect 4593 7349 4595 7383
rect 4747 7349 4749 7383
rect 4749 7349 4781 7383
rect 4819 7349 4851 7383
rect 4851 7349 4853 7383
rect 5005 7349 5007 7383
rect 5007 7349 5039 7383
rect 5077 7349 5109 7383
rect 5109 7349 5111 7383
rect 5263 7349 5265 7383
rect 5265 7349 5297 7383
rect 5335 7349 5367 7383
rect 5367 7349 5369 7383
rect 5521 7349 5523 7383
rect 5523 7349 5555 7383
rect 5593 7349 5625 7383
rect 5625 7349 5627 7383
rect 5779 7349 5781 7383
rect 5781 7349 5813 7383
rect 5851 7349 5883 7383
rect 5883 7349 5885 7383
rect 6037 7349 6039 7383
rect 6039 7349 6071 7383
rect 6109 7349 6141 7383
rect 6141 7349 6143 7383
rect 3622 7262 3656 7264
rect 3622 7230 3656 7262
rect 3622 7160 3656 7192
rect 3622 7158 3656 7160
rect 3880 7262 3914 7264
rect 3880 7230 3914 7262
rect 3880 7160 3914 7192
rect 3880 7158 3914 7160
rect 4138 7262 4172 7264
rect 4138 7230 4172 7262
rect 4138 7160 4172 7192
rect 4138 7158 4172 7160
rect 4396 7262 4430 7264
rect 4396 7230 4430 7262
rect 4396 7160 4430 7192
rect 4396 7158 4430 7160
rect 4654 7262 4688 7264
rect 4654 7230 4688 7262
rect 4654 7160 4688 7192
rect 4654 7158 4688 7160
rect 4912 7262 4946 7264
rect 4912 7230 4946 7262
rect 4912 7160 4946 7192
rect 4912 7158 4946 7160
rect 5170 7262 5204 7264
rect 5170 7230 5204 7262
rect 5170 7160 5204 7192
rect 5170 7158 5204 7160
rect 5428 7262 5462 7264
rect 5428 7230 5462 7262
rect 5428 7160 5462 7192
rect 5428 7158 5462 7160
rect 5686 7262 5720 7264
rect 5686 7230 5720 7262
rect 5686 7160 5720 7192
rect 5686 7158 5720 7160
rect 5944 7262 5978 7264
rect 5944 7230 5978 7262
rect 5944 7160 5978 7192
rect 5944 7158 5978 7160
rect 6202 7262 6236 7264
rect 6202 7230 6236 7262
rect 6202 7160 6236 7192
rect 6202 7158 6236 7160
rect 3715 7039 3717 7073
rect 3717 7039 3749 7073
rect 3787 7039 3819 7073
rect 3819 7039 3821 7073
rect 6037 7039 6039 7073
rect 6039 7039 6071 7073
rect 6109 7039 6141 7073
rect 6141 7039 6143 7073
rect 3715 6931 3717 6965
rect 3717 6931 3749 6965
rect 3787 6931 3819 6965
rect 3819 6931 3821 6965
rect 3973 6931 3975 6965
rect 3975 6931 4007 6965
rect 4045 6931 4077 6965
rect 4077 6931 4079 6965
rect 4231 6931 4233 6965
rect 4233 6931 4265 6965
rect 4303 6931 4335 6965
rect 4335 6931 4337 6965
rect 5005 6931 5007 6965
rect 5007 6931 5039 6965
rect 5077 6931 5109 6965
rect 5109 6931 5111 6965
rect 5263 6931 5265 6965
rect 5265 6931 5297 6965
rect 5335 6931 5367 6965
rect 5367 6931 5369 6965
rect 6037 6931 6039 6965
rect 6039 6931 6071 6965
rect 6109 6931 6141 6965
rect 6141 6931 6143 6965
rect 3622 6844 3656 6846
rect 3622 6812 3656 6844
rect 3622 6742 3656 6774
rect 3622 6740 3656 6742
rect 3880 6844 3914 6846
rect 3880 6812 3914 6844
rect 3880 6742 3914 6774
rect 3880 6740 3914 6742
rect 4138 6844 4172 6846
rect 4138 6812 4172 6844
rect 4138 6742 4172 6774
rect 4138 6740 4172 6742
rect 4396 6844 4430 6846
rect 4396 6812 4430 6844
rect 4396 6742 4430 6774
rect 4396 6740 4430 6742
rect 4654 6844 4688 6846
rect 4654 6812 4688 6844
rect 4654 6742 4688 6774
rect 4654 6740 4688 6742
rect 4912 6844 4946 6846
rect 4912 6812 4946 6844
rect 4912 6742 4946 6774
rect 4912 6740 4946 6742
rect 5170 6844 5204 6846
rect 5170 6812 5204 6844
rect 5170 6742 5204 6774
rect 5170 6740 5204 6742
rect 5428 6844 5462 6846
rect 5428 6812 5462 6844
rect 5428 6742 5462 6774
rect 5428 6740 5462 6742
rect 5686 6844 5720 6846
rect 5686 6812 5720 6844
rect 5686 6742 5720 6774
rect 5686 6740 5720 6742
rect 5944 6844 5978 6846
rect 5944 6812 5978 6844
rect 5944 6742 5978 6774
rect 5944 6740 5978 6742
rect 6202 6844 6236 6846
rect 6202 6812 6236 6844
rect 6202 6742 6236 6774
rect 6202 6740 6236 6742
rect 3715 6621 3717 6655
rect 3717 6621 3749 6655
rect 3787 6621 3819 6655
rect 3819 6621 3821 6655
rect 4489 6621 4491 6655
rect 4491 6621 4523 6655
rect 4561 6621 4593 6655
rect 4593 6621 4595 6655
rect 4747 6621 4749 6655
rect 4749 6621 4781 6655
rect 4819 6621 4851 6655
rect 4851 6621 4853 6655
rect 5521 6621 5523 6655
rect 5523 6621 5555 6655
rect 5593 6621 5625 6655
rect 5625 6621 5627 6655
rect 5779 6621 5781 6655
rect 5781 6621 5813 6655
rect 5851 6621 5883 6655
rect 5883 6621 5885 6655
rect 6037 6621 6039 6655
rect 6039 6621 6071 6655
rect 6109 6621 6141 6655
rect 6141 6621 6143 6655
rect 3715 6513 3717 6547
rect 3717 6513 3749 6547
rect 3787 6513 3819 6547
rect 3819 6513 3821 6547
rect 4489 6513 4491 6547
rect 4491 6513 4523 6547
rect 4561 6513 4593 6547
rect 4593 6513 4595 6547
rect 4747 6513 4749 6547
rect 4749 6513 4781 6547
rect 4819 6513 4851 6547
rect 4851 6513 4853 6547
rect 5521 6513 5523 6547
rect 5523 6513 5555 6547
rect 5593 6513 5625 6547
rect 5625 6513 5627 6547
rect 5779 6513 5781 6547
rect 5781 6513 5813 6547
rect 5851 6513 5883 6547
rect 5883 6513 5885 6547
rect 6037 6513 6039 6547
rect 6039 6513 6071 6547
rect 6109 6513 6141 6547
rect 6141 6513 6143 6547
rect 3622 6426 3656 6428
rect 3622 6394 3656 6426
rect 3622 6324 3656 6356
rect 3622 6322 3656 6324
rect 3880 6426 3914 6428
rect 3880 6394 3914 6426
rect 3880 6324 3914 6356
rect 3880 6322 3914 6324
rect 4138 6426 4172 6428
rect 4138 6394 4172 6426
rect 4138 6324 4172 6356
rect 4138 6322 4172 6324
rect 4396 6426 4430 6428
rect 4396 6394 4430 6426
rect 4396 6324 4430 6356
rect 4396 6322 4430 6324
rect 4654 6426 4688 6428
rect 4654 6394 4688 6426
rect 4654 6324 4688 6356
rect 4654 6322 4688 6324
rect 4912 6426 4946 6428
rect 4912 6394 4946 6426
rect 4912 6324 4946 6356
rect 4912 6322 4946 6324
rect 5170 6426 5204 6428
rect 5170 6394 5204 6426
rect 5170 6324 5204 6356
rect 5170 6322 5204 6324
rect 5428 6426 5462 6428
rect 5428 6394 5462 6426
rect 5428 6324 5462 6356
rect 5428 6322 5462 6324
rect 5686 6426 5720 6428
rect 5686 6394 5720 6426
rect 5686 6324 5720 6356
rect 5686 6322 5720 6324
rect 5944 6426 5978 6428
rect 5944 6394 5978 6426
rect 5944 6324 5978 6356
rect 5944 6322 5978 6324
rect 6202 6426 6236 6428
rect 6202 6394 6236 6426
rect 6202 6324 6236 6356
rect 6202 6322 6236 6324
rect 3715 6203 3717 6237
rect 3717 6203 3749 6237
rect 3787 6203 3819 6237
rect 3819 6203 3821 6237
rect 3973 6203 3975 6237
rect 3975 6203 4007 6237
rect 4045 6203 4077 6237
rect 4077 6203 4079 6237
rect 4231 6203 4233 6237
rect 4233 6203 4265 6237
rect 4303 6203 4335 6237
rect 4335 6203 4337 6237
rect 5005 6203 5007 6237
rect 5007 6203 5039 6237
rect 5077 6203 5109 6237
rect 5109 6203 5111 6237
rect 5263 6203 5265 6237
rect 5265 6203 5297 6237
rect 5335 6203 5367 6237
rect 5367 6203 5369 6237
rect 6037 6203 6039 6237
rect 6039 6203 6071 6237
rect 6109 6203 6141 6237
rect 6141 6203 6143 6237
rect 3715 6095 3717 6129
rect 3717 6095 3749 6129
rect 3787 6095 3819 6129
rect 3819 6095 3821 6129
rect 3973 6095 3975 6129
rect 3975 6095 4007 6129
rect 4045 6095 4077 6129
rect 4077 6095 4079 6129
rect 4231 6095 4233 6129
rect 4233 6095 4265 6129
rect 4303 6095 4335 6129
rect 4335 6095 4337 6129
rect 5005 6095 5007 6129
rect 5007 6095 5039 6129
rect 5077 6095 5109 6129
rect 5109 6095 5111 6129
rect 5263 6095 5265 6129
rect 5265 6095 5297 6129
rect 5335 6095 5367 6129
rect 5367 6095 5369 6129
rect 6037 6095 6039 6129
rect 6039 6095 6071 6129
rect 6109 6095 6141 6129
rect 6141 6095 6143 6129
rect 3622 6008 3656 6010
rect 3622 5976 3656 6008
rect 3622 5906 3656 5938
rect 3622 5904 3656 5906
rect 3880 6008 3914 6010
rect 3880 5976 3914 6008
rect 3880 5906 3914 5938
rect 3880 5904 3914 5906
rect 4138 6008 4172 6010
rect 4138 5976 4172 6008
rect 4138 5906 4172 5938
rect 4138 5904 4172 5906
rect 4396 6008 4430 6010
rect 4396 5976 4430 6008
rect 4396 5906 4430 5938
rect 4396 5904 4430 5906
rect 4654 6008 4688 6010
rect 4654 5976 4688 6008
rect 4654 5906 4688 5938
rect 4654 5904 4688 5906
rect 4912 6008 4946 6010
rect 4912 5976 4946 6008
rect 4912 5906 4946 5938
rect 4912 5904 4946 5906
rect 5170 6008 5204 6010
rect 5170 5976 5204 6008
rect 5170 5906 5204 5938
rect 5170 5904 5204 5906
rect 5428 6008 5462 6010
rect 5428 5976 5462 6008
rect 5428 5906 5462 5938
rect 5428 5904 5462 5906
rect 5686 6008 5720 6010
rect 5686 5976 5720 6008
rect 5686 5906 5720 5938
rect 5686 5904 5720 5906
rect 5944 6008 5978 6010
rect 5944 5976 5978 6008
rect 5944 5906 5978 5938
rect 5944 5904 5978 5906
rect 6202 6008 6236 6010
rect 6202 5976 6236 6008
rect 6202 5906 6236 5938
rect 6202 5904 6236 5906
rect 3715 5785 3717 5819
rect 3717 5785 3749 5819
rect 3787 5785 3819 5819
rect 3819 5785 3821 5819
rect 4489 5785 4491 5819
rect 4491 5785 4523 5819
rect 4561 5785 4593 5819
rect 4593 5785 4595 5819
rect 4747 5785 4749 5819
rect 4749 5785 4781 5819
rect 4819 5785 4851 5819
rect 4851 5785 4853 5819
rect 5521 5785 5523 5819
rect 5523 5785 5555 5819
rect 5593 5785 5625 5819
rect 5625 5785 5627 5819
rect 5779 5785 5781 5819
rect 5781 5785 5813 5819
rect 5851 5785 5883 5819
rect 5883 5785 5885 5819
rect 6037 5785 6039 5819
rect 6039 5785 6071 5819
rect 6109 5785 6141 5819
rect 6141 5785 6143 5819
rect 3715 5677 3717 5711
rect 3717 5677 3749 5711
rect 3787 5677 3819 5711
rect 3819 5677 3821 5711
rect 4489 5677 4491 5711
rect 4491 5677 4523 5711
rect 4561 5677 4593 5711
rect 4593 5677 4595 5711
rect 4747 5677 4749 5711
rect 4749 5677 4781 5711
rect 4819 5677 4851 5711
rect 4851 5677 4853 5711
rect 5521 5677 5523 5711
rect 5523 5677 5555 5711
rect 5593 5677 5625 5711
rect 5625 5677 5627 5711
rect 5779 5677 5781 5711
rect 5781 5677 5813 5711
rect 5851 5677 5883 5711
rect 5883 5677 5885 5711
rect 6037 5677 6039 5711
rect 6039 5677 6071 5711
rect 6109 5677 6141 5711
rect 6141 5677 6143 5711
rect 3622 5590 3656 5592
rect 3622 5558 3656 5590
rect 3622 5488 3656 5520
rect 3622 5486 3656 5488
rect 3880 5590 3914 5592
rect 3880 5558 3914 5590
rect 3880 5488 3914 5520
rect 3880 5486 3914 5488
rect 4138 5590 4172 5592
rect 4138 5558 4172 5590
rect 4138 5488 4172 5520
rect 4138 5486 4172 5488
rect 4396 5590 4430 5592
rect 4396 5558 4430 5590
rect 4396 5488 4430 5520
rect 4396 5486 4430 5488
rect 4654 5590 4688 5592
rect 4654 5558 4688 5590
rect 4654 5488 4688 5520
rect 4654 5486 4688 5488
rect 4912 5590 4946 5592
rect 4912 5558 4946 5590
rect 4912 5488 4946 5520
rect 4912 5486 4946 5488
rect 5170 5590 5204 5592
rect 5170 5558 5204 5590
rect 5170 5488 5204 5520
rect 5170 5486 5204 5488
rect 5428 5590 5462 5592
rect 5428 5558 5462 5590
rect 5428 5488 5462 5520
rect 5428 5486 5462 5488
rect 5686 5590 5720 5592
rect 5686 5558 5720 5590
rect 5686 5488 5720 5520
rect 5686 5486 5720 5488
rect 5944 5590 5978 5592
rect 5944 5558 5978 5590
rect 5944 5488 5978 5520
rect 5944 5486 5978 5488
rect 6202 5590 6236 5592
rect 6202 5558 6236 5590
rect 6202 5488 6236 5520
rect 6202 5486 6236 5488
rect 3715 5367 3717 5401
rect 3717 5367 3749 5401
rect 3787 5367 3819 5401
rect 3819 5367 3821 5401
rect 3973 5367 3975 5401
rect 3975 5367 4007 5401
rect 4045 5367 4077 5401
rect 4077 5367 4079 5401
rect 4231 5367 4233 5401
rect 4233 5367 4265 5401
rect 4303 5367 4335 5401
rect 4335 5367 4337 5401
rect 5005 5367 5007 5401
rect 5007 5367 5039 5401
rect 5077 5367 5109 5401
rect 5109 5367 5111 5401
rect 5263 5367 5265 5401
rect 5265 5367 5297 5401
rect 5335 5367 5367 5401
rect 5367 5367 5369 5401
rect 6037 5367 6039 5401
rect 6039 5367 6071 5401
rect 6109 5367 6141 5401
rect 6141 5367 6143 5401
rect 3715 5259 3717 5293
rect 3717 5259 3749 5293
rect 3787 5259 3819 5293
rect 3819 5259 3821 5293
rect 3973 5259 3975 5293
rect 3975 5259 4007 5293
rect 4045 5259 4077 5293
rect 4077 5259 4079 5293
rect 4231 5259 4233 5293
rect 4233 5259 4265 5293
rect 4303 5259 4335 5293
rect 4335 5259 4337 5293
rect 5005 5259 5007 5293
rect 5007 5259 5039 5293
rect 5077 5259 5109 5293
rect 5109 5259 5111 5293
rect 5263 5259 5265 5293
rect 5265 5259 5297 5293
rect 5335 5259 5367 5293
rect 5367 5259 5369 5293
rect 6037 5259 6039 5293
rect 6039 5259 6071 5293
rect 6109 5259 6141 5293
rect 6141 5259 6143 5293
rect 3622 5172 3656 5174
rect 3622 5140 3656 5172
rect 3622 5070 3656 5102
rect 3622 5068 3656 5070
rect 3880 5172 3914 5174
rect 3880 5140 3914 5172
rect 3880 5070 3914 5102
rect 3880 5068 3914 5070
rect 4138 5172 4172 5174
rect 4138 5140 4172 5172
rect 4138 5070 4172 5102
rect 4138 5068 4172 5070
rect 4396 5172 4430 5174
rect 4396 5140 4430 5172
rect 4396 5070 4430 5102
rect 4396 5068 4430 5070
rect 4654 5172 4688 5174
rect 4654 5140 4688 5172
rect 4654 5070 4688 5102
rect 4654 5068 4688 5070
rect 4912 5172 4946 5174
rect 4912 5140 4946 5172
rect 4912 5070 4946 5102
rect 4912 5068 4946 5070
rect 5170 5172 5204 5174
rect 5170 5140 5204 5172
rect 5170 5070 5204 5102
rect 5170 5068 5204 5070
rect 5428 5172 5462 5174
rect 5428 5140 5462 5172
rect 5428 5070 5462 5102
rect 5428 5068 5462 5070
rect 5686 5172 5720 5174
rect 5686 5140 5720 5172
rect 5686 5070 5720 5102
rect 5686 5068 5720 5070
rect 5944 5172 5978 5174
rect 5944 5140 5978 5172
rect 5944 5070 5978 5102
rect 5944 5068 5978 5070
rect 6202 5172 6236 5174
rect 6202 5140 6236 5172
rect 6202 5070 6236 5102
rect 6202 5068 6236 5070
rect 3715 4949 3717 4983
rect 3717 4949 3749 4983
rect 3787 4949 3819 4983
rect 3819 4949 3821 4983
rect 4489 4949 4491 4983
rect 4491 4949 4523 4983
rect 4561 4949 4593 4983
rect 4593 4949 4595 4983
rect 4747 4949 4749 4983
rect 4749 4949 4781 4983
rect 4819 4949 4851 4983
rect 4851 4949 4853 4983
rect 5521 4949 5523 4983
rect 5523 4949 5555 4983
rect 5593 4949 5625 4983
rect 5625 4949 5627 4983
rect 5779 4949 5781 4983
rect 5781 4949 5813 4983
rect 5851 4949 5883 4983
rect 5883 4949 5885 4983
rect 6037 4949 6039 4983
rect 6039 4949 6071 4983
rect 6109 4949 6141 4983
rect 6141 4949 6143 4983
rect 3715 4841 3717 4875
rect 3717 4841 3749 4875
rect 3787 4841 3819 4875
rect 3819 4841 3821 4875
rect 4489 4841 4491 4875
rect 4491 4841 4523 4875
rect 4561 4841 4593 4875
rect 4593 4841 4595 4875
rect 4747 4841 4749 4875
rect 4749 4841 4781 4875
rect 4819 4841 4851 4875
rect 4851 4841 4853 4875
rect 5521 4841 5523 4875
rect 5523 4841 5555 4875
rect 5593 4841 5625 4875
rect 5625 4841 5627 4875
rect 5779 4841 5781 4875
rect 5781 4841 5813 4875
rect 5851 4841 5883 4875
rect 5883 4841 5885 4875
rect 6037 4841 6039 4875
rect 6039 4841 6071 4875
rect 6109 4841 6141 4875
rect 6141 4841 6143 4875
rect 3622 4754 3656 4756
rect 3622 4722 3656 4754
rect 3622 4652 3656 4684
rect 3622 4650 3656 4652
rect 3880 4754 3914 4756
rect 3880 4722 3914 4754
rect 3880 4652 3914 4684
rect 3880 4650 3914 4652
rect 4138 4754 4172 4756
rect 4138 4722 4172 4754
rect 4138 4652 4172 4684
rect 4138 4650 4172 4652
rect 4396 4754 4430 4756
rect 4396 4722 4430 4754
rect 4396 4652 4430 4684
rect 4396 4650 4430 4652
rect 4654 4754 4688 4756
rect 4654 4722 4688 4754
rect 4654 4652 4688 4684
rect 4654 4650 4688 4652
rect 4912 4754 4946 4756
rect 4912 4722 4946 4754
rect 4912 4652 4946 4684
rect 4912 4650 4946 4652
rect 5170 4754 5204 4756
rect 5170 4722 5204 4754
rect 5170 4652 5204 4684
rect 5170 4650 5204 4652
rect 5428 4754 5462 4756
rect 5428 4722 5462 4754
rect 5428 4652 5462 4684
rect 5428 4650 5462 4652
rect 5686 4754 5720 4756
rect 5686 4722 5720 4754
rect 5686 4652 5720 4684
rect 5686 4650 5720 4652
rect 5944 4754 5978 4756
rect 5944 4722 5978 4754
rect 5944 4652 5978 4684
rect 5944 4650 5978 4652
rect 6202 4754 6236 4756
rect 6202 4722 6236 4754
rect 6202 4652 6236 4684
rect 6202 4650 6236 4652
rect 3715 4531 3717 4565
rect 3717 4531 3749 4565
rect 3787 4531 3819 4565
rect 3819 4531 3821 4565
rect 3973 4531 3975 4565
rect 3975 4531 4007 4565
rect 4045 4531 4077 4565
rect 4077 4531 4079 4565
rect 4231 4531 4233 4565
rect 4233 4531 4265 4565
rect 4303 4531 4335 4565
rect 4335 4531 4337 4565
rect 5005 4531 5007 4565
rect 5007 4531 5039 4565
rect 5077 4531 5109 4565
rect 5109 4531 5111 4565
rect 5263 4531 5265 4565
rect 5265 4531 5297 4565
rect 5335 4531 5367 4565
rect 5367 4531 5369 4565
rect 6037 4531 6039 4565
rect 6039 4531 6071 4565
rect 6109 4531 6141 4565
rect 6141 4531 6143 4565
rect 3715 4423 3717 4457
rect 3717 4423 3749 4457
rect 3787 4423 3819 4457
rect 3819 4423 3821 4457
rect 3973 4423 3975 4457
rect 3975 4423 4007 4457
rect 4045 4423 4077 4457
rect 4077 4423 4079 4457
rect 4231 4423 4233 4457
rect 4233 4423 4265 4457
rect 4303 4423 4335 4457
rect 4335 4423 4337 4457
rect 4489 4423 4491 4457
rect 4491 4423 4523 4457
rect 4561 4423 4593 4457
rect 4593 4423 4595 4457
rect 4747 4423 4749 4457
rect 4749 4423 4781 4457
rect 4819 4423 4851 4457
rect 4851 4423 4853 4457
rect 5005 4423 5007 4457
rect 5007 4423 5039 4457
rect 5077 4423 5109 4457
rect 5109 4423 5111 4457
rect 5263 4423 5265 4457
rect 5265 4423 5297 4457
rect 5335 4423 5367 4457
rect 5367 4423 5369 4457
rect 5521 4423 5523 4457
rect 5523 4423 5555 4457
rect 5593 4423 5625 4457
rect 5625 4423 5627 4457
rect 5779 4423 5781 4457
rect 5781 4423 5813 4457
rect 5851 4423 5883 4457
rect 5883 4423 5885 4457
rect 6037 4423 6039 4457
rect 6039 4423 6071 4457
rect 6109 4423 6141 4457
rect 6141 4423 6143 4457
rect 3622 4336 3656 4338
rect 3622 4304 3656 4336
rect 3622 4234 3656 4266
rect 3622 4232 3656 4234
rect 3880 4336 3914 4338
rect 3880 4304 3914 4336
rect 3880 4234 3914 4266
rect 3880 4232 3914 4234
rect 4138 4336 4172 4338
rect 4138 4304 4172 4336
rect 4138 4234 4172 4266
rect 4138 4232 4172 4234
rect 4396 4336 4430 4338
rect 4396 4304 4430 4336
rect 4396 4234 4430 4266
rect 4396 4232 4430 4234
rect 4654 4336 4688 4338
rect 4654 4304 4688 4336
rect 4654 4234 4688 4266
rect 4654 4232 4688 4234
rect 4912 4336 4946 4338
rect 4912 4304 4946 4336
rect 4912 4234 4946 4266
rect 4912 4232 4946 4234
rect 5170 4336 5204 4338
rect 5170 4304 5204 4336
rect 5170 4234 5204 4266
rect 5170 4232 5204 4234
rect 5428 4336 5462 4338
rect 5428 4304 5462 4336
rect 5428 4234 5462 4266
rect 5428 4232 5462 4234
rect 5686 4336 5720 4338
rect 5686 4304 5720 4336
rect 5686 4234 5720 4266
rect 5686 4232 5720 4234
rect 5944 4336 5978 4338
rect 5944 4304 5978 4336
rect 5944 4234 5978 4266
rect 5944 4232 5978 4234
rect 6202 4336 6236 4338
rect 6202 4304 6236 4336
rect 6202 4234 6236 4266
rect 6202 4232 6236 4234
rect 6316 4235 6350 4238
rect 6316 4204 6350 4235
rect 3715 4113 3717 4147
rect 3717 4113 3749 4147
rect 3787 4113 3819 4147
rect 3819 4113 3821 4147
rect 6037 4113 6039 4147
rect 6039 4113 6071 4147
rect 6109 4113 6141 4147
rect 6141 4113 6143 4147
rect 8451 6938 8453 6972
rect 8453 6938 8485 6972
rect 8523 6938 8555 6972
rect 8555 6938 8557 6972
rect 8709 6938 8711 6972
rect 8711 6938 8743 6972
rect 8781 6938 8813 6972
rect 8813 6938 8815 6972
rect 8967 6938 8969 6972
rect 8969 6938 9001 6972
rect 9039 6938 9071 6972
rect 9071 6938 9073 6972
rect 9225 6938 9227 6972
rect 9227 6938 9259 6972
rect 9297 6938 9329 6972
rect 9329 6938 9331 6972
rect 9483 6938 9485 6972
rect 9485 6938 9517 6972
rect 9555 6938 9587 6972
rect 9587 6938 9589 6972
rect 9741 6938 9743 6972
rect 9743 6938 9775 6972
rect 9813 6938 9845 6972
rect 9845 6938 9847 6972
rect 8358 6851 8392 6853
rect 8358 6819 8392 6851
rect 8358 6749 8392 6781
rect 8358 6747 8392 6749
rect 8616 6851 8650 6853
rect 8616 6819 8650 6851
rect 8616 6749 8650 6781
rect 8616 6747 8650 6749
rect 8874 6851 8908 6853
rect 8874 6819 8908 6851
rect 8874 6749 8908 6781
rect 8874 6747 8908 6749
rect 9132 6851 9166 6853
rect 9132 6819 9166 6851
rect 9132 6749 9166 6781
rect 9132 6747 9166 6749
rect 9390 6851 9424 6853
rect 9390 6819 9424 6851
rect 9390 6749 9424 6781
rect 9390 6747 9424 6749
rect 9648 6851 9682 6853
rect 9648 6819 9682 6851
rect 9648 6749 9682 6781
rect 9648 6747 9682 6749
rect 9906 6851 9940 6853
rect 9906 6819 9940 6851
rect 9906 6749 9940 6781
rect 9906 6747 9940 6749
rect 8451 6628 8453 6662
rect 8453 6628 8485 6662
rect 8523 6628 8555 6662
rect 8555 6628 8557 6662
rect 9741 6628 9743 6662
rect 9743 6628 9775 6662
rect 9813 6628 9845 6662
rect 9845 6628 9847 6662
rect 8451 6520 8453 6554
rect 8453 6520 8485 6554
rect 8523 6520 8555 6554
rect 8555 6520 8557 6554
rect 8709 6520 8711 6554
rect 8711 6520 8743 6554
rect 8781 6520 8813 6554
rect 8813 6520 8815 6554
rect 8967 6520 8969 6554
rect 8969 6520 9001 6554
rect 9039 6520 9071 6554
rect 9071 6520 9073 6554
rect 9225 6520 9227 6554
rect 9227 6520 9259 6554
rect 9297 6520 9329 6554
rect 9329 6520 9331 6554
rect 9483 6520 9485 6554
rect 9485 6520 9517 6554
rect 9555 6520 9587 6554
rect 9587 6520 9589 6554
rect 9741 6520 9743 6554
rect 9743 6520 9775 6554
rect 9813 6520 9845 6554
rect 9845 6520 9847 6554
rect 8358 6433 8392 6435
rect 8358 6401 8392 6433
rect 8358 6331 8392 6363
rect 8358 6329 8392 6331
rect 8616 6433 8650 6435
rect 8616 6401 8650 6433
rect 8616 6331 8650 6363
rect 8616 6329 8650 6331
rect 8874 6433 8908 6435
rect 8874 6401 8908 6433
rect 8874 6331 8908 6363
rect 8874 6329 8908 6331
rect 9132 6433 9166 6435
rect 9132 6401 9166 6433
rect 9132 6331 9166 6363
rect 9132 6329 9166 6331
rect 9390 6433 9424 6435
rect 9390 6401 9424 6433
rect 9390 6331 9424 6363
rect 9390 6329 9424 6331
rect 9648 6433 9682 6435
rect 9648 6401 9682 6433
rect 9648 6331 9682 6363
rect 9648 6329 9682 6331
rect 9906 6433 9940 6435
rect 9906 6401 9940 6433
rect 9906 6331 9940 6363
rect 9906 6329 9940 6331
rect 8451 6210 8453 6244
rect 8453 6210 8485 6244
rect 8523 6210 8555 6244
rect 8555 6210 8557 6244
rect 9741 6210 9743 6244
rect 9743 6210 9775 6244
rect 9813 6210 9845 6244
rect 9845 6210 9847 6244
rect 8451 6102 8453 6136
rect 8453 6102 8485 6136
rect 8523 6102 8555 6136
rect 8555 6102 8557 6136
rect 8709 6102 8711 6136
rect 8711 6102 8743 6136
rect 8781 6102 8813 6136
rect 8813 6102 8815 6136
rect 8967 6102 8969 6136
rect 8969 6102 9001 6136
rect 9039 6102 9071 6136
rect 9071 6102 9073 6136
rect 9225 6102 9227 6136
rect 9227 6102 9259 6136
rect 9297 6102 9329 6136
rect 9329 6102 9331 6136
rect 9483 6102 9485 6136
rect 9485 6102 9517 6136
rect 9555 6102 9587 6136
rect 9587 6102 9589 6136
rect 9741 6102 9743 6136
rect 9743 6102 9775 6136
rect 9813 6102 9845 6136
rect 9845 6102 9847 6136
rect 8358 6015 8392 6017
rect 8358 5983 8392 6015
rect 8358 5913 8392 5945
rect 8358 5911 8392 5913
rect 8616 6015 8650 6017
rect 8616 5983 8650 6015
rect 8616 5913 8650 5945
rect 8616 5911 8650 5913
rect 8874 6015 8908 6017
rect 8874 5983 8908 6015
rect 8874 5913 8908 5945
rect 8874 5911 8908 5913
rect 9132 6015 9166 6017
rect 9132 5983 9166 6015
rect 9132 5913 9166 5945
rect 9132 5911 9166 5913
rect 9390 6015 9424 6017
rect 9390 5983 9424 6015
rect 9390 5913 9424 5945
rect 9390 5911 9424 5913
rect 9648 6015 9682 6017
rect 9648 5983 9682 6015
rect 9648 5913 9682 5945
rect 9648 5911 9682 5913
rect 9906 6015 9940 6017
rect 9906 5983 9940 6015
rect 9906 5913 9940 5945
rect 9906 5911 9940 5913
rect 8451 5792 8453 5826
rect 8453 5792 8485 5826
rect 8523 5792 8555 5826
rect 8555 5792 8557 5826
rect 9741 5792 9743 5826
rect 9743 5792 9775 5826
rect 9813 5792 9845 5826
rect 9845 5792 9847 5826
rect 8451 5684 8453 5718
rect 8453 5684 8485 5718
rect 8523 5684 8555 5718
rect 8555 5684 8557 5718
rect 8709 5684 8711 5718
rect 8711 5684 8743 5718
rect 8781 5684 8813 5718
rect 8813 5684 8815 5718
rect 8967 5684 8969 5718
rect 8969 5684 9001 5718
rect 9039 5684 9071 5718
rect 9071 5684 9073 5718
rect 9225 5684 9227 5718
rect 9227 5684 9259 5718
rect 9297 5684 9329 5718
rect 9329 5684 9331 5718
rect 9483 5684 9485 5718
rect 9485 5684 9517 5718
rect 9555 5684 9587 5718
rect 9587 5684 9589 5718
rect 9741 5684 9743 5718
rect 9743 5684 9775 5718
rect 9813 5684 9845 5718
rect 9845 5684 9847 5718
rect 8358 5597 8392 5599
rect 8358 5565 8392 5597
rect 8358 5495 8392 5527
rect 8358 5493 8392 5495
rect 8616 5597 8650 5599
rect 8616 5565 8650 5597
rect 8616 5495 8650 5527
rect 8616 5493 8650 5495
rect 8874 5597 8908 5599
rect 8874 5565 8908 5597
rect 8874 5495 8908 5527
rect 8874 5493 8908 5495
rect 9132 5597 9166 5599
rect 9132 5565 9166 5597
rect 9132 5495 9166 5527
rect 9132 5493 9166 5495
rect 9390 5597 9424 5599
rect 9390 5565 9424 5597
rect 9390 5495 9424 5527
rect 9390 5493 9424 5495
rect 9648 5597 9682 5599
rect 9648 5565 9682 5597
rect 9648 5495 9682 5527
rect 9648 5493 9682 5495
rect 9906 5597 9940 5599
rect 9906 5565 9940 5597
rect 9906 5495 9940 5527
rect 9906 5493 9940 5495
rect 8451 5374 8453 5408
rect 8453 5374 8485 5408
rect 8523 5374 8555 5408
rect 8555 5374 8557 5408
rect 9741 5374 9743 5408
rect 9743 5374 9775 5408
rect 9813 5374 9845 5408
rect 9845 5374 9847 5408
rect 8451 5266 8453 5300
rect 8453 5266 8485 5300
rect 8523 5266 8555 5300
rect 8555 5266 8557 5300
rect 8709 5266 8711 5300
rect 8711 5266 8743 5300
rect 8781 5266 8813 5300
rect 8813 5266 8815 5300
rect 8967 5266 8969 5300
rect 8969 5266 9001 5300
rect 9039 5266 9071 5300
rect 9071 5266 9073 5300
rect 9225 5266 9227 5300
rect 9227 5266 9259 5300
rect 9297 5266 9329 5300
rect 9329 5266 9331 5300
rect 9483 5266 9485 5300
rect 9485 5266 9517 5300
rect 9555 5266 9587 5300
rect 9587 5266 9589 5300
rect 9741 5266 9743 5300
rect 9743 5266 9775 5300
rect 9813 5266 9845 5300
rect 9845 5266 9847 5300
rect 8358 5179 8392 5181
rect 8358 5147 8392 5179
rect 8358 5077 8392 5109
rect 8358 5075 8392 5077
rect 8616 5179 8650 5181
rect 8616 5147 8650 5179
rect 8616 5077 8650 5109
rect 8616 5075 8650 5077
rect 8874 5179 8908 5181
rect 8874 5147 8908 5179
rect 8874 5077 8908 5109
rect 8874 5075 8908 5077
rect 9132 5179 9166 5181
rect 9132 5147 9166 5179
rect 9132 5077 9166 5109
rect 9132 5075 9166 5077
rect 9390 5179 9424 5181
rect 9390 5147 9424 5179
rect 9390 5077 9424 5109
rect 9390 5075 9424 5077
rect 9648 5179 9682 5181
rect 9648 5147 9682 5179
rect 9648 5077 9682 5109
rect 9648 5075 9682 5077
rect 9906 5179 9940 5181
rect 9906 5147 9940 5179
rect 9906 5077 9940 5109
rect 9906 5075 9940 5077
rect 8451 4956 8453 4990
rect 8453 4956 8485 4990
rect 8523 4956 8555 4990
rect 8555 4956 8557 4990
rect 9741 4956 9743 4990
rect 9743 4956 9775 4990
rect 9813 4956 9845 4990
rect 9845 4956 9847 4990
rect 8451 4848 8453 4882
rect 8453 4848 8485 4882
rect 8523 4848 8555 4882
rect 8555 4848 8557 4882
rect 8709 4848 8711 4882
rect 8711 4848 8743 4882
rect 8781 4848 8813 4882
rect 8813 4848 8815 4882
rect 8967 4848 8969 4882
rect 8969 4848 9001 4882
rect 9039 4848 9071 4882
rect 9071 4848 9073 4882
rect 9225 4848 9227 4882
rect 9227 4848 9259 4882
rect 9297 4848 9329 4882
rect 9329 4848 9331 4882
rect 9483 4848 9485 4882
rect 9485 4848 9517 4882
rect 9555 4848 9587 4882
rect 9587 4848 9589 4882
rect 9741 4848 9743 4882
rect 9743 4848 9775 4882
rect 9813 4848 9845 4882
rect 9845 4848 9847 4882
rect 8358 4761 8392 4763
rect 8358 4729 8392 4761
rect 8358 4659 8392 4691
rect 8358 4657 8392 4659
rect 8616 4761 8650 4763
rect 8616 4729 8650 4761
rect 8616 4659 8650 4691
rect 8616 4657 8650 4659
rect 8874 4761 8908 4763
rect 8874 4729 8908 4761
rect 8874 4659 8908 4691
rect 8874 4657 8908 4659
rect 9132 4761 9166 4763
rect 9132 4729 9166 4761
rect 9132 4659 9166 4691
rect 9132 4657 9166 4659
rect 9390 4761 9424 4763
rect 9390 4729 9424 4761
rect 9390 4659 9424 4691
rect 9390 4657 9424 4659
rect 9648 4761 9682 4763
rect 9648 4729 9682 4761
rect 9648 4659 9682 4691
rect 9648 4657 9682 4659
rect 9906 4761 9940 4763
rect 9906 4729 9940 4761
rect 9906 4659 9940 4691
rect 9906 4657 9940 4659
rect 8451 4538 8453 4572
rect 8453 4538 8485 4572
rect 8523 4538 8555 4572
rect 8555 4538 8557 4572
rect 9741 4538 9743 4572
rect 9743 4538 9775 4572
rect 9813 4538 9845 4572
rect 9845 4538 9847 4572
rect 8451 4430 8453 4464
rect 8453 4430 8485 4464
rect 8523 4430 8555 4464
rect 8555 4430 8557 4464
rect 8709 4430 8711 4464
rect 8711 4430 8743 4464
rect 8781 4430 8813 4464
rect 8813 4430 8815 4464
rect 8967 4430 8969 4464
rect 8969 4430 9001 4464
rect 9039 4430 9071 4464
rect 9071 4430 9073 4464
rect 9225 4430 9227 4464
rect 9227 4430 9259 4464
rect 9297 4430 9329 4464
rect 9329 4430 9331 4464
rect 9483 4430 9485 4464
rect 9485 4430 9517 4464
rect 9555 4430 9587 4464
rect 9587 4430 9589 4464
rect 9741 4430 9743 4464
rect 9743 4430 9775 4464
rect 9813 4430 9845 4464
rect 9845 4430 9847 4464
rect 8358 4343 8392 4345
rect 8358 4311 8392 4343
rect 8358 4241 8392 4273
rect 8358 4239 8392 4241
rect 8616 4343 8650 4345
rect 8616 4311 8650 4343
rect 8616 4241 8650 4273
rect 8616 4239 8650 4241
rect 8874 4343 8908 4345
rect 8874 4311 8908 4343
rect 8874 4241 8908 4273
rect 8874 4239 8908 4241
rect 9132 4343 9166 4345
rect 9132 4311 9166 4343
rect 9132 4241 9166 4273
rect 9132 4239 9166 4241
rect 9390 4343 9424 4345
rect 9390 4311 9424 4343
rect 9390 4241 9424 4273
rect 9390 4239 9424 4241
rect 9648 4343 9682 4345
rect 9648 4311 9682 4343
rect 9648 4241 9682 4273
rect 9648 4239 9682 4241
rect 9906 4343 9940 4345
rect 9906 4311 9940 4343
rect 9906 4241 9940 4273
rect 9906 4239 9940 4241
rect 8451 4120 8453 4154
rect 8453 4120 8485 4154
rect 8523 4120 8555 4154
rect 8555 4120 8557 4154
rect 9741 4120 9743 4154
rect 9743 4120 9775 4154
rect 9813 4120 9845 4154
rect 9845 4120 9847 4154
rect 9906 4018 9940 4052
rect -2115 3916 -2113 3950
rect -2113 3916 -2081 3950
rect -2043 3916 -2011 3950
rect -2011 3916 -2009 3950
rect 1239 3916 1241 3950
rect 1241 3916 1273 3950
rect 1311 3916 1343 3950
rect 1343 3916 1345 3950
<< metal1 >>
rect -945 11213 12450 11259
rect -945 10892 -899 11213
rect 3077 10913 5187 10959
rect -1245 10846 766 10892
rect -1245 10663 -1199 10846
rect -1245 10629 -1239 10663
rect -1205 10629 -1199 10663
rect -1245 10567 -1199 10629
rect -987 10567 -941 10846
rect -1245 10561 -941 10567
rect -1245 10527 -1146 10561
rect -1112 10527 -1074 10561
rect -1040 10527 -941 10561
rect -1245 10521 -941 10527
rect -1245 10433 -1199 10521
rect -1245 10399 -1239 10433
rect -1205 10399 -1199 10433
rect -1245 10361 -1199 10399
rect -1245 10327 -1239 10361
rect -1205 10327 -1199 10361
rect -1245 10239 -1199 10327
rect -987 10433 -941 10521
rect -987 10399 -981 10433
rect -947 10399 -941 10433
rect -987 10361 -941 10399
rect -987 10327 -981 10361
rect -947 10327 -941 10361
rect -987 10239 -941 10327
rect -732 10433 -680 10480
rect -732 10399 -723 10433
rect -689 10399 -680 10433
rect -732 10361 -680 10399
rect -732 10327 -723 10361
rect -689 10327 -680 10361
rect -732 10242 -680 10327
rect -471 10433 -425 10846
rect 45 10567 91 10846
rect 303 10567 349 10846
rect 45 10561 349 10567
rect 45 10527 144 10561
rect 178 10527 216 10561
rect 250 10527 349 10561
rect 45 10521 349 10527
rect -471 10399 -465 10433
rect -431 10399 -425 10433
rect -471 10361 -425 10399
rect -471 10327 -465 10361
rect -431 10327 -425 10361
rect -1245 10233 -941 10239
rect -1245 10199 -1146 10233
rect -1112 10199 -1074 10233
rect -1040 10199 -941 10233
rect -1245 10193 -941 10199
rect -1245 10131 -1199 10193
rect -987 10131 -941 10193
rect -913 10190 -897 10242
rect -845 10190 -825 10242
rect -773 10190 -639 10242
rect -587 10190 -567 10242
rect -515 10190 -499 10242
rect -1245 10125 -941 10131
rect -1245 10091 -1146 10125
rect -1112 10091 -1074 10125
rect -1040 10091 -941 10125
rect -1245 10085 -941 10091
rect -1245 9997 -1199 10085
rect -1245 9963 -1239 9997
rect -1205 9963 -1199 9997
rect -1245 9925 -1199 9963
rect -1245 9891 -1239 9925
rect -1205 9891 -1199 9925
rect -1245 9803 -1199 9891
rect -987 9997 -941 10085
rect -913 10082 -897 10134
rect -845 10082 -825 10134
rect -773 10082 -757 10134
rect -655 10082 -639 10134
rect -587 10082 -567 10134
rect -515 10082 -499 10134
rect -987 9963 -981 9997
rect -947 9963 -941 9997
rect -987 9925 -941 9963
rect -987 9891 -981 9925
rect -947 9891 -941 9925
rect -987 9803 -941 9891
rect -732 10006 -680 10044
rect -732 9934 -680 9954
rect -732 9844 -680 9882
rect -471 9997 -425 10327
rect -216 10442 -164 10480
rect -216 10370 -164 10390
rect -216 10280 -164 10318
rect 45 10433 91 10521
rect 45 10399 51 10433
rect 85 10399 91 10433
rect 45 10361 91 10399
rect 45 10327 51 10361
rect 85 10327 91 10361
rect -397 10190 -381 10242
rect -329 10190 -309 10242
rect -257 10190 -241 10242
rect -139 10190 -123 10242
rect -71 10190 -51 10242
rect 1 10190 17 10242
rect 45 10239 91 10327
rect 303 10433 349 10521
rect 303 10399 309 10433
rect 343 10399 349 10433
rect 303 10361 349 10399
rect 303 10327 309 10361
rect 343 10327 349 10361
rect 303 10239 349 10327
rect 45 10233 349 10239
rect 45 10199 144 10233
rect 178 10199 216 10233
rect 250 10199 349 10233
rect 45 10193 349 10199
rect -397 10082 -381 10134
rect -329 10082 -309 10134
rect -257 10082 -123 10134
rect -71 10082 -51 10134
rect 1 10082 17 10134
rect 45 10131 91 10193
rect 303 10131 349 10193
rect 45 10125 349 10131
rect 45 10091 144 10125
rect 178 10091 216 10125
rect 250 10091 349 10125
rect 45 10085 349 10091
rect -471 9963 -465 9997
rect -431 9963 -425 9997
rect -471 9925 -425 9963
rect -471 9891 -465 9925
rect -431 9891 -425 9925
rect -1245 9797 -941 9803
rect -1245 9763 -1146 9797
rect -1112 9763 -1074 9797
rect -1040 9763 -941 9797
rect -1245 9757 -941 9763
rect -1245 9695 -1199 9757
rect -987 9695 -941 9757
rect -1245 9689 -941 9695
rect -1245 9655 -1146 9689
rect -1112 9655 -1074 9689
rect -1040 9655 -941 9689
rect -1245 9649 -941 9655
rect -1245 9561 -1199 9649
rect -1245 9527 -1239 9561
rect -1205 9527 -1199 9561
rect -1245 9489 -1199 9527
rect -1245 9455 -1239 9489
rect -1205 9455 -1199 9489
rect -1245 9367 -1199 9455
rect -987 9561 -941 9649
rect -987 9527 -981 9561
rect -947 9527 -941 9561
rect -987 9489 -941 9527
rect -987 9455 -981 9489
rect -947 9455 -941 9489
rect -987 9367 -941 9455
rect -732 9561 -680 9608
rect -732 9527 -723 9561
rect -689 9527 -680 9561
rect -732 9489 -680 9527
rect -732 9455 -723 9489
rect -689 9455 -680 9489
rect -732 9370 -680 9455
rect -471 9561 -425 9891
rect -216 9997 -164 10082
rect -216 9963 -207 9997
rect -173 9963 -164 9997
rect -216 9925 -164 9963
rect -216 9891 -207 9925
rect -173 9891 -164 9925
rect -216 9844 -164 9891
rect 45 9997 91 10085
rect 45 9963 51 9997
rect 85 9963 91 9997
rect 45 9925 91 9963
rect 45 9891 51 9925
rect 85 9891 91 9925
rect 45 9803 91 9891
rect 303 9997 349 10085
rect 303 9963 309 9997
rect 343 9963 349 9997
rect 303 9925 349 9963
rect 303 9891 309 9925
rect 343 9891 349 9925
rect 303 9803 349 9891
rect 45 9797 349 9803
rect 45 9763 144 9797
rect 178 9763 216 9797
rect 250 9763 349 9797
rect 45 9757 349 9763
rect 45 9695 91 9757
rect 303 9695 349 9757
rect 45 9689 349 9695
rect 45 9655 144 9689
rect 178 9655 216 9689
rect 250 9655 349 9689
rect 45 9649 349 9655
rect -471 9527 -465 9561
rect -431 9527 -425 9561
rect -471 9489 -425 9527
rect -471 9455 -465 9489
rect -431 9455 -425 9489
rect -1245 9361 -941 9367
rect -1245 9327 -1146 9361
rect -1112 9327 -1074 9361
rect -1040 9327 -941 9361
rect -1245 9321 -941 9327
rect -1245 9259 -1199 9321
rect -987 9259 -941 9321
rect -913 9318 -897 9370
rect -845 9318 -825 9370
rect -773 9318 -639 9370
rect -587 9318 -567 9370
rect -515 9318 -499 9370
rect -1245 9253 -941 9259
rect -1245 9219 -1146 9253
rect -1112 9219 -1074 9253
rect -1040 9219 -941 9253
rect -1245 9213 -941 9219
rect -1245 9125 -1199 9213
rect -1245 9091 -1239 9125
rect -1205 9091 -1199 9125
rect -1245 9053 -1199 9091
rect -1245 9019 -1239 9053
rect -1205 9019 -1199 9053
rect -1245 8931 -1199 9019
rect -987 9125 -941 9213
rect -913 9210 -897 9262
rect -845 9210 -825 9262
rect -773 9210 -757 9262
rect -655 9210 -639 9262
rect -587 9210 -567 9262
rect -515 9210 -499 9262
rect -987 9091 -981 9125
rect -947 9091 -941 9125
rect -987 9053 -941 9091
rect -987 9019 -981 9053
rect -947 9019 -941 9053
rect -987 8931 -941 9019
rect -732 9134 -680 9172
rect -732 9062 -680 9082
rect -732 8972 -680 9010
rect -471 9125 -425 9455
rect -216 9570 -164 9608
rect -216 9498 -164 9518
rect -216 9408 -164 9446
rect 45 9561 91 9649
rect 45 9527 51 9561
rect 85 9527 91 9561
rect 45 9489 91 9527
rect 45 9455 51 9489
rect 85 9455 91 9489
rect -397 9318 -381 9370
rect -329 9318 -309 9370
rect -257 9318 -241 9370
rect -139 9318 -123 9370
rect -71 9318 -51 9370
rect 1 9318 17 9370
rect 45 9367 91 9455
rect 303 9561 349 9649
rect 303 9527 309 9561
rect 343 9527 349 9561
rect 303 9489 349 9527
rect 303 9455 309 9489
rect 343 9455 349 9489
rect 303 9367 349 9455
rect 45 9361 349 9367
rect 45 9327 144 9361
rect 178 9327 216 9361
rect 250 9327 349 9361
rect 45 9321 349 9327
rect -397 9210 -381 9262
rect -329 9210 -309 9262
rect -257 9210 -123 9262
rect -71 9210 -51 9262
rect 1 9210 17 9262
rect 45 9259 91 9321
rect 303 9259 349 9321
rect 45 9253 349 9259
rect 45 9219 144 9253
rect 178 9219 216 9253
rect 250 9219 349 9253
rect 45 9213 349 9219
rect -471 9091 -465 9125
rect -431 9091 -425 9125
rect -471 9053 -425 9091
rect -471 9019 -465 9053
rect -431 9019 -425 9053
rect -1245 8925 -941 8931
rect -1245 8891 -1146 8925
rect -1112 8891 -1074 8925
rect -1040 8891 -941 8925
rect -1245 8885 -941 8891
rect -471 8875 -425 9019
rect -216 9125 -164 9210
rect -216 9091 -207 9125
rect -173 9091 -164 9125
rect -216 9053 -164 9091
rect -216 9019 -207 9053
rect -173 9019 -164 9053
rect -216 8972 -164 9019
rect 45 9125 91 9213
rect 45 9091 51 9125
rect 85 9091 91 9125
rect 45 9053 91 9091
rect 45 9019 51 9053
rect 85 9019 91 9053
rect 45 8931 91 9019
rect 303 9125 349 9213
rect 303 9091 309 9125
rect 343 9091 349 9125
rect 303 9053 349 9091
rect 303 9019 309 9053
rect 343 9019 349 9053
rect 303 8931 349 9019
rect 45 8925 349 8931
rect 45 8891 144 8925
rect 178 8891 216 8925
rect 250 8891 349 8925
rect 45 8885 349 8891
rect 3077 10777 3123 10913
rect 3077 10771 3593 10777
rect 3077 10737 3176 10771
rect 3210 10737 3248 10771
rect 3282 10737 3434 10771
rect 3468 10737 3506 10771
rect 3540 10737 3593 10771
rect 3077 10731 3593 10737
rect 3077 10652 3123 10731
rect 3077 10618 3083 10652
rect 3117 10618 3123 10652
rect 3077 10580 3123 10618
rect 3077 10546 3083 10580
rect 3117 10546 3123 10580
rect 3077 10467 3123 10546
rect 3335 10652 3381 10731
rect 3649 10728 3683 10780
rect 3735 10728 3755 10780
rect 3807 10728 3841 10780
rect 4423 10728 4457 10780
rect 4509 10728 4529 10780
rect 4581 10728 4615 10780
rect 5141 10777 5187 10913
rect 4671 10771 5187 10777
rect 4671 10737 4724 10771
rect 4758 10737 4796 10771
rect 4830 10737 4982 10771
rect 5016 10737 5054 10771
rect 5088 10737 5187 10771
rect 4671 10731 5187 10737
rect 3335 10618 3341 10652
rect 3375 10618 3381 10652
rect 3335 10580 3381 10618
rect 3335 10546 3341 10580
rect 3375 10546 3381 10580
rect 3335 10499 3381 10546
rect 3590 10661 3642 10699
rect 3590 10589 3642 10609
rect 3590 10499 3642 10537
rect 3851 10652 3897 10699
rect 3851 10618 3857 10652
rect 3891 10618 3897 10652
rect 3851 10580 3897 10618
rect 3851 10546 3857 10580
rect 3891 10546 3897 10580
rect 3077 10461 3307 10467
rect 3077 10427 3176 10461
rect 3210 10427 3248 10461
rect 3282 10427 3307 10461
rect 3077 10421 3307 10427
rect 3077 10359 3123 10421
rect 3077 10353 3307 10359
rect 3077 10319 3176 10353
rect 3210 10319 3248 10353
rect 3282 10319 3307 10353
rect 3077 10313 3307 10319
rect 3077 10234 3123 10313
rect 3077 10200 3083 10234
rect 3117 10200 3123 10234
rect 3077 10162 3123 10200
rect 3077 10128 3083 10162
rect 3117 10128 3123 10162
rect 3077 10049 3123 10128
rect 3335 10234 3381 10357
rect 3335 10200 3341 10234
rect 3375 10200 3381 10234
rect 3335 10162 3381 10200
rect 3335 10128 3341 10162
rect 3375 10128 3381 10162
rect 3077 10043 3307 10049
rect 3077 10009 3176 10043
rect 3210 10009 3248 10043
rect 3282 10009 3307 10043
rect 3077 10003 3307 10009
rect 3077 9941 3123 10003
rect 3077 9935 3307 9941
rect 3077 9901 3176 9935
rect 3210 9901 3248 9935
rect 3282 9901 3307 9935
rect 3077 9895 3307 9901
rect 3077 9816 3123 9895
rect 3077 9782 3083 9816
rect 3117 9782 3123 9816
rect 3077 9744 3123 9782
rect 3077 9710 3083 9744
rect 3117 9710 3123 9744
rect 3077 9631 3123 9710
rect 3335 9816 3381 10128
rect 3590 10243 3642 10281
rect 3590 10171 3642 10191
rect 3590 10081 3642 10119
rect 3851 10234 3897 10546
rect 4106 10661 4158 10699
rect 4106 10589 4158 10609
rect 4106 10499 4158 10537
rect 4367 10652 4413 10699
rect 4367 10618 4373 10652
rect 4407 10618 4413 10652
rect 4367 10580 4413 10618
rect 4367 10546 4373 10580
rect 4407 10546 4413 10580
rect 3925 10415 3941 10467
rect 3993 10415 4013 10467
rect 4065 10415 4099 10467
rect 4165 10415 4199 10467
rect 4251 10415 4271 10467
rect 4323 10415 4339 10467
rect 3925 10310 3941 10362
rect 3993 10310 4013 10362
rect 4065 10310 4099 10362
rect 4165 10310 4199 10362
rect 4251 10310 4271 10362
rect 4323 10310 4339 10362
rect 3851 10200 3857 10234
rect 3891 10200 3897 10234
rect 3851 10162 3897 10200
rect 3851 10128 3857 10162
rect 3891 10128 3897 10162
rect 3409 9997 3425 10049
rect 3477 9997 3497 10049
rect 3549 9997 3583 10049
rect 3649 9997 3683 10049
rect 3735 9997 3755 10049
rect 3807 9997 3823 10049
rect 3409 9892 3425 9944
rect 3477 9892 3497 9944
rect 3549 9892 3583 9944
rect 3649 9892 3683 9944
rect 3735 9892 3755 9944
rect 3807 9892 3823 9944
rect 3335 9782 3341 9816
rect 3375 9782 3381 9816
rect 3335 9744 3381 9782
rect 3335 9710 3341 9744
rect 3375 9710 3381 9744
rect 3077 9625 3307 9631
rect 3077 9591 3176 9625
rect 3210 9591 3248 9625
rect 3282 9591 3307 9625
rect 3077 9585 3307 9591
rect 3077 9523 3123 9585
rect 3077 9517 3307 9523
rect 3077 9483 3176 9517
rect 3210 9483 3248 9517
rect 3282 9483 3307 9517
rect 3077 9477 3307 9483
rect 3077 9398 3123 9477
rect 3077 9364 3083 9398
rect 3117 9364 3123 9398
rect 3077 9326 3123 9364
rect 3077 9292 3083 9326
rect 3117 9292 3123 9326
rect 3077 9213 3123 9292
rect 3335 9398 3381 9710
rect 3590 9825 3642 9863
rect 3590 9753 3642 9773
rect 3590 9663 3642 9701
rect 3851 9816 3897 10128
rect 4106 10243 4158 10281
rect 4106 10171 4158 10191
rect 4106 10081 4158 10119
rect 4367 10234 4413 10546
rect 4622 10661 4674 10699
rect 4622 10589 4674 10609
rect 4622 10499 4674 10537
rect 4883 10652 4929 10731
rect 4883 10618 4889 10652
rect 4923 10618 4929 10652
rect 4883 10580 4929 10618
rect 4883 10546 4889 10580
rect 4923 10546 4929 10580
rect 4883 10499 4929 10546
rect 5141 10652 5187 10731
rect 5141 10618 5147 10652
rect 5181 10618 5187 10652
rect 5141 10580 5187 10618
rect 5141 10546 5147 10580
rect 5181 10546 5187 10580
rect 5141 10464 5187 10546
rect 4957 10458 5187 10464
rect 4957 10424 4982 10458
rect 5016 10424 5054 10458
rect 5088 10424 5187 10458
rect 4957 10418 5187 10424
rect 4367 10200 4373 10234
rect 4407 10200 4413 10234
rect 4367 10162 4413 10200
rect 4367 10128 4373 10162
rect 4407 10128 4413 10162
rect 3851 9782 3857 9816
rect 3891 9782 3897 9816
rect 3851 9744 3897 9782
rect 3851 9710 3857 9744
rect 3891 9710 3897 9744
rect 3335 9364 3341 9398
rect 3375 9364 3381 9398
rect 3335 9326 3381 9364
rect 3335 9292 3341 9326
rect 3375 9292 3381 9326
rect 3077 9207 3307 9213
rect 3077 9173 3176 9207
rect 3210 9173 3248 9207
rect 3282 9173 3307 9207
rect 3077 9167 3307 9173
rect 3077 9101 3123 9167
rect 3077 9095 3307 9101
rect 3077 9061 3176 9095
rect 3210 9061 3248 9095
rect 3282 9061 3307 9095
rect 3077 9055 3307 9061
rect 3077 8976 3123 9055
rect 3077 8942 3083 8976
rect 3117 8942 3123 8976
rect 3077 8904 3123 8942
rect 3077 8870 3083 8904
rect 3117 8870 3123 8904
rect 3077 8791 3123 8870
rect 3335 8976 3381 9292
rect 3590 9407 3642 9445
rect 3590 9335 3642 9355
rect 3590 9245 3642 9283
rect 3851 9398 3897 9710
rect 4106 9825 4158 9863
rect 4106 9753 4158 9773
rect 4106 9663 4158 9701
rect 4367 9816 4413 10128
rect 4622 10243 4674 10281
rect 4622 10171 4674 10191
rect 4622 10081 4674 10119
rect 4883 10234 4929 10370
rect 5141 10359 5187 10418
rect 4957 10353 5187 10359
rect 4957 10319 4982 10353
rect 5016 10319 5054 10353
rect 5088 10319 5187 10353
rect 4957 10313 5187 10319
rect 4883 10200 4889 10234
rect 4923 10200 4929 10234
rect 4883 10162 4929 10200
rect 4883 10128 4889 10162
rect 4923 10128 4929 10162
rect 4441 9997 4457 10049
rect 4509 9997 4529 10049
rect 4581 9997 4615 10049
rect 4681 9997 4715 10049
rect 4767 9997 4787 10049
rect 4839 9997 4855 10049
rect 4441 9892 4457 9944
rect 4509 9892 4529 9944
rect 4581 9892 4615 9944
rect 4681 9892 4715 9944
rect 4767 9892 4787 9944
rect 4839 9892 4855 9944
rect 4367 9782 4373 9816
rect 4407 9782 4413 9816
rect 4367 9744 4413 9782
rect 4367 9710 4373 9744
rect 4407 9710 4413 9744
rect 3925 9579 3941 9631
rect 3993 9579 4013 9631
rect 4065 9579 4099 9631
rect 4165 9579 4199 9631
rect 4251 9579 4271 9631
rect 4323 9579 4339 9631
rect 3925 9474 3941 9526
rect 3993 9474 4013 9526
rect 4065 9474 4099 9526
rect 4165 9474 4199 9526
rect 4251 9474 4271 9526
rect 4323 9474 4339 9526
rect 3851 9364 3857 9398
rect 3891 9364 3897 9398
rect 3851 9326 3897 9364
rect 3851 9292 3857 9326
rect 3891 9292 3897 9326
rect 3409 9161 3425 9213
rect 3477 9161 3497 9213
rect 3549 9161 3583 9213
rect 3649 9161 3683 9213
rect 3735 9161 3755 9213
rect 3807 9161 3823 9213
rect 3409 9052 3425 9104
rect 3477 9052 3497 9104
rect 3549 9052 3583 9104
rect 3649 9052 3683 9104
rect 3735 9052 3755 9104
rect 3807 9052 3823 9104
rect 3335 8942 3341 8976
rect 3375 8942 3381 8976
rect 3335 8904 3381 8942
rect 3335 8870 3341 8904
rect 3375 8870 3381 8904
rect 3077 8785 3307 8791
rect 3077 8751 3176 8785
rect 3210 8751 3248 8785
rect 3282 8751 3307 8785
rect 3077 8745 3307 8751
rect 3335 8781 3381 8870
rect 3590 8985 3642 9023
rect 3590 8913 3642 8933
rect 3590 8823 3642 8861
rect 3851 8976 3897 9292
rect 4106 9407 4158 9445
rect 4106 9335 4158 9355
rect 4106 9245 4158 9283
rect 4367 9398 4413 9710
rect 4622 9825 4674 9863
rect 4622 9753 4674 9773
rect 4622 9663 4674 9701
rect 4883 9816 4929 10128
rect 5141 10234 5187 10313
rect 5141 10200 5147 10234
rect 5181 10200 5187 10234
rect 5141 10162 5187 10200
rect 5141 10128 5147 10162
rect 5181 10128 5187 10162
rect 5141 10049 5187 10128
rect 4957 10043 5187 10049
rect 4957 10009 4982 10043
rect 5016 10009 5054 10043
rect 5088 10009 5187 10043
rect 4957 10003 5187 10009
rect 5141 9941 5187 10003
rect 4957 9935 5187 9941
rect 4957 9901 4982 9935
rect 5016 9901 5054 9935
rect 5088 9901 5187 9935
rect 4957 9895 5187 9901
rect 4883 9782 4889 9816
rect 4923 9782 4929 9816
rect 4883 9744 4929 9782
rect 4883 9710 4889 9744
rect 4923 9710 4929 9744
rect 4367 9364 4373 9398
rect 4407 9364 4413 9398
rect 4367 9326 4413 9364
rect 4367 9292 4373 9326
rect 4407 9292 4413 9326
rect 3851 8942 3857 8976
rect 3891 8942 3897 8976
rect 3851 8904 3897 8942
rect 3851 8870 3857 8904
rect 3891 8870 3897 8904
rect 3851 8781 3897 8870
rect 4106 8985 4158 9023
rect 4106 8913 4158 8933
rect 4106 8823 4158 8861
rect 4367 8976 4413 9292
rect 4622 9407 4674 9445
rect 4622 9335 4674 9355
rect 4622 9245 4674 9283
rect 4883 9398 4929 9710
rect 5141 9816 5187 9895
rect 5141 9782 5147 9816
rect 5181 9782 5187 9816
rect 5141 9744 5187 9782
rect 5141 9710 5147 9744
rect 5181 9710 5187 9744
rect 5141 9628 5187 9710
rect 4957 9622 5187 9628
rect 4957 9588 4982 9622
rect 5016 9588 5054 9622
rect 5088 9588 5187 9622
rect 4957 9582 5187 9588
rect 5141 9523 5187 9582
rect 4957 9517 5187 9523
rect 4957 9483 4982 9517
rect 5016 9483 5054 9517
rect 5088 9483 5187 9517
rect 4957 9477 5187 9483
rect 4883 9364 4889 9398
rect 4923 9364 4929 9398
rect 4883 9326 4929 9364
rect 4883 9292 4889 9326
rect 4923 9292 4929 9326
rect 4441 9161 4457 9213
rect 4509 9161 4529 9213
rect 4581 9161 4615 9213
rect 4681 9161 4715 9213
rect 4767 9161 4787 9213
rect 4839 9161 4855 9213
rect 4441 9052 4457 9104
rect 4509 9052 4529 9104
rect 4581 9052 4615 9104
rect 4681 9052 4715 9104
rect 4767 9052 4787 9104
rect 4839 9052 4855 9104
rect 4367 8942 4373 8976
rect 4407 8942 4413 8976
rect 4367 8904 4413 8942
rect 4367 8870 4373 8904
rect 4407 8870 4413 8904
rect 3077 8679 3123 8745
rect 3335 8735 3897 8781
rect 3925 8739 3941 8791
rect 3993 8739 4013 8791
rect 4065 8739 4099 8791
rect 4165 8739 4199 8791
rect 4251 8739 4271 8791
rect 4323 8739 4339 8791
rect 4367 8781 4413 8870
rect 4622 8985 4674 9023
rect 4622 8913 4674 8933
rect 4622 8823 4674 8861
rect 4883 8976 4929 9292
rect 5141 9398 5187 9477
rect 5141 9364 5147 9398
rect 5181 9364 5187 9398
rect 5141 9326 5187 9364
rect 5141 9292 5147 9326
rect 5181 9292 5187 9326
rect 5141 9210 5187 9292
rect 4957 9204 5187 9210
rect 4957 9170 4982 9204
rect 5016 9170 5054 9204
rect 5088 9170 5187 9204
rect 4957 9164 5187 9170
rect 5141 9101 5187 9164
rect 4957 9095 5187 9101
rect 4957 9061 4982 9095
rect 5016 9061 5054 9095
rect 5088 9061 5187 9095
rect 4957 9055 5187 9061
rect 4883 8942 4889 8976
rect 4923 8942 4929 8976
rect 4883 8904 4929 8942
rect 4883 8870 4889 8904
rect 4923 8870 4929 8904
rect 4883 8781 4929 8870
rect 5141 8976 5187 9055
rect 5141 8942 5147 8976
rect 5181 8942 5187 8976
rect 5141 8904 5187 8942
rect 5141 8870 5147 8904
rect 5181 8870 5187 8904
rect 5141 8788 5187 8870
rect 3077 8673 3307 8679
rect 3077 8639 3176 8673
rect 3210 8639 3248 8673
rect 3282 8639 3307 8673
rect 3077 8633 3307 8639
rect 3077 8554 3123 8633
rect 3077 8520 3083 8554
rect 3117 8520 3123 8554
rect 3077 8482 3123 8520
rect 3077 8448 3083 8482
rect 3117 8448 3123 8482
rect 2227 8371 2307 8383
rect 2227 8319 2241 8371
rect 2293 8369 2307 8371
rect 3077 8369 3123 8448
rect 3335 8554 3381 8601
rect 3335 8520 3341 8554
rect 3375 8520 3381 8554
rect 3335 8482 3381 8520
rect 3335 8448 3341 8482
rect 3375 8448 3381 8482
rect 3335 8369 3381 8448
rect 3590 8563 3642 8601
rect 3590 8491 3642 8511
rect 3590 8401 3642 8439
rect 3851 8554 3897 8735
rect 4367 8735 4929 8781
rect 4957 8782 5187 8788
rect 4957 8748 4982 8782
rect 5016 8748 5054 8782
rect 5088 8748 5187 8782
rect 4957 8742 5187 8748
rect 3925 8630 3941 8682
rect 3993 8630 4013 8682
rect 4065 8630 4099 8682
rect 4165 8630 4199 8682
rect 4251 8630 4271 8682
rect 4323 8630 4339 8682
rect 3851 8520 3857 8554
rect 3891 8520 3897 8554
rect 3851 8482 3897 8520
rect 3851 8448 3857 8482
rect 3891 8448 3897 8482
rect 2293 8363 3593 8369
rect 2293 8329 2969 8363
rect 3003 8329 3176 8363
rect 3210 8329 3248 8363
rect 3282 8329 3434 8363
rect 3468 8329 3506 8363
rect 3540 8329 3593 8363
rect 2293 8323 3593 8329
rect 2293 8319 2307 8323
rect 2227 8307 2307 8319
rect 3649 8317 3683 8369
rect 3735 8317 3755 8369
rect 3807 8317 3823 8369
rect -2214 8186 1444 8232
rect -2214 8028 -2168 8186
rect -1956 8031 -1910 8186
rect -1701 8031 -1649 8186
rect -1440 8031 -1394 8186
rect -1185 8031 -1133 8186
rect 879 8031 931 8186
rect 1140 8031 1186 8186
rect -1956 8028 -924 8031
rect -2214 8022 -924 8028
rect -2214 7988 -2115 8022
rect -2081 7988 -2043 8022
rect -2009 7988 -1857 8022
rect -1823 7988 -1785 8022
rect -1751 7988 -1599 8022
rect -1565 7988 -1527 8022
rect -1493 7988 -1341 8022
rect -1307 7988 -1269 8022
rect -1235 7988 -1083 8022
rect -1049 7988 -1011 8022
rect -977 7988 -924 8022
rect -2214 7982 -924 7988
rect -2214 7903 -2168 7982
rect -2214 7869 -2208 7903
rect -2174 7869 -2168 7903
rect -2214 7831 -2168 7869
rect -2214 7797 -2208 7831
rect -2174 7797 -2168 7831
rect -2214 7718 -2168 7797
rect -1956 7979 -924 7982
rect -850 7979 -834 8031
rect -782 7979 -762 8031
rect -710 7979 -676 8031
rect -610 7979 -576 8031
rect -524 7979 -504 8031
rect -452 7979 -436 8031
rect -334 7979 -318 8031
rect -266 7979 -246 8031
rect -194 7979 -160 8031
rect -94 7979 -60 8031
rect -8 7979 12 8031
rect 64 7979 80 8031
rect 182 7979 198 8031
rect 250 7979 270 8031
rect 322 7979 356 8031
rect 422 7979 456 8031
rect 508 7979 528 8031
rect 580 7979 596 8031
rect 670 8028 1186 8031
rect 1398 8028 1444 8186
rect 670 8022 1444 8028
rect 670 7988 723 8022
rect 757 7988 795 8022
rect 829 7988 981 8022
rect 1015 7988 1053 8022
rect 1087 7988 1239 8022
rect 1273 7988 1311 8022
rect 1345 7988 1444 8022
rect 670 7982 1444 7988
rect 3851 7982 3897 8448
rect 4106 8563 4158 8601
rect 4106 8491 4158 8511
rect 4106 8401 4158 8439
rect 4367 8554 4413 8735
rect 5141 8679 5187 8742
rect 4957 8673 5187 8679
rect 4957 8639 4982 8673
rect 5016 8639 5054 8673
rect 5088 8639 5187 8673
rect 4957 8633 5187 8639
rect 4367 8520 4373 8554
rect 4407 8520 4413 8554
rect 4367 8482 4413 8520
rect 4367 8448 4373 8482
rect 4407 8448 4413 8482
rect 4367 7982 4413 8448
rect 4622 8563 4674 8601
rect 4622 8491 4674 8511
rect 4622 8401 4674 8439
rect 4883 8554 4929 8601
rect 4883 8520 4889 8554
rect 4923 8520 4929 8554
rect 4883 8482 4929 8520
rect 4883 8448 4889 8482
rect 4923 8448 4929 8482
rect 4883 8369 4929 8448
rect 5141 8554 5187 8633
rect 5141 8520 5147 8554
rect 5181 8520 5187 8554
rect 5141 8482 5187 8520
rect 5141 8448 5147 8482
rect 5181 8448 5187 8482
rect 5141 8369 5187 8448
rect 4441 8317 4457 8369
rect 4509 8317 4529 8369
rect 4581 8317 4615 8369
rect 4671 8363 5187 8369
rect 4671 8329 4724 8363
rect 4758 8329 4796 8363
rect 4830 8329 4982 8363
rect 5016 8329 5054 8363
rect 5088 8329 5187 8363
rect 4671 8323 5187 8329
rect 7003 10885 7049 11213
rect 7261 10885 7307 11213
rect 7003 10879 7307 10885
rect 7003 10845 7102 10879
rect 7136 10845 7174 10879
rect 7208 10845 7307 10879
rect 7003 10839 7307 10845
rect 7003 10751 7049 10839
rect 7003 10717 7009 10751
rect 7043 10717 7049 10751
rect 7003 10679 7049 10717
rect 7003 10645 7009 10679
rect 7043 10645 7049 10679
rect 7003 10557 7049 10645
rect 7261 10751 7307 10839
rect 7261 10717 7267 10751
rect 7301 10717 7307 10751
rect 7261 10679 7307 10717
rect 7261 10645 7267 10679
rect 7301 10645 7307 10679
rect 7261 10557 7307 10645
rect 7519 10751 7565 10885
rect 7519 10717 7525 10751
rect 7559 10717 7565 10751
rect 7519 10679 7565 10717
rect 7519 10645 7525 10679
rect 7559 10645 7565 10679
rect 7003 10551 7307 10557
rect 7003 10517 7102 10551
rect 7136 10517 7174 10551
rect 7208 10517 7307 10551
rect 7003 10511 7307 10517
rect 7003 10449 7049 10511
rect 7261 10449 7307 10511
rect 7335 10508 7351 10560
rect 7403 10508 7423 10560
rect 7475 10508 7491 10560
rect 7003 10443 7307 10449
rect 7003 10409 7102 10443
rect 7136 10409 7174 10443
rect 7208 10409 7307 10443
rect 7003 10403 7307 10409
rect 7003 10315 7049 10403
rect 7003 10281 7009 10315
rect 7043 10281 7049 10315
rect 7003 10243 7049 10281
rect 7003 10209 7009 10243
rect 7043 10209 7049 10243
rect 7003 10121 7049 10209
rect 7261 10315 7307 10403
rect 7335 10400 7351 10452
rect 7403 10400 7423 10452
rect 7475 10400 7491 10452
rect 7261 10281 7267 10315
rect 7301 10281 7307 10315
rect 7261 10243 7307 10281
rect 7261 10209 7267 10243
rect 7301 10209 7307 10243
rect 7261 10121 7307 10209
rect 7003 10115 7307 10121
rect 7003 10081 7102 10115
rect 7136 10081 7174 10115
rect 7208 10081 7307 10115
rect 7003 10075 7307 10081
rect 7003 10013 7049 10075
rect 7261 10013 7307 10075
rect 7003 10007 7307 10013
rect 7003 9973 7102 10007
rect 7136 9973 7174 10007
rect 7208 9973 7307 10007
rect 7003 9967 7307 9973
rect 7003 9879 7049 9967
rect 7003 9845 7009 9879
rect 7043 9845 7049 9879
rect 7003 9807 7049 9845
rect 7003 9773 7009 9807
rect 7043 9773 7049 9807
rect 7003 9685 7049 9773
rect 7261 9879 7307 9967
rect 7261 9845 7267 9879
rect 7301 9845 7307 9879
rect 7261 9807 7307 9845
rect 7261 9773 7267 9807
rect 7301 9773 7307 9807
rect 7261 9685 7307 9773
rect 7519 10315 7565 10645
rect 7777 10751 7823 11213
rect 8293 10981 8339 11213
rect 8293 10947 8299 10981
rect 8333 10947 8339 10981
rect 8293 10885 8339 10947
rect 8551 10885 8597 11213
rect 7777 10717 7783 10751
rect 7817 10717 7823 10751
rect 7777 10679 7823 10717
rect 7777 10645 7783 10679
rect 7817 10645 7823 10679
rect 7593 10508 7609 10560
rect 7661 10508 7681 10560
rect 7733 10508 7749 10560
rect 7593 10400 7609 10452
rect 7661 10400 7681 10452
rect 7733 10400 7749 10452
rect 7519 10281 7525 10315
rect 7559 10281 7565 10315
rect 7519 10243 7565 10281
rect 7519 10209 7525 10243
rect 7559 10209 7565 10243
rect 7519 9879 7565 10209
rect 7519 9845 7525 9879
rect 7559 9845 7565 9879
rect 7519 9807 7565 9845
rect 7519 9773 7525 9807
rect 7559 9773 7565 9807
rect 7003 9679 7307 9685
rect 7003 9645 7102 9679
rect 7136 9645 7174 9679
rect 7208 9645 7307 9679
rect 7003 9639 7307 9645
rect 7003 9577 7049 9639
rect 7261 9577 7307 9639
rect 7335 9636 7351 9688
rect 7403 9636 7423 9688
rect 7475 9636 7491 9688
rect 7003 9571 7307 9577
rect 7003 9537 7102 9571
rect 7136 9537 7174 9571
rect 7208 9537 7307 9571
rect 7003 9531 7307 9537
rect 7003 9443 7049 9531
rect 7003 9409 7009 9443
rect 7043 9409 7049 9443
rect 7003 9371 7049 9409
rect 7003 9337 7009 9371
rect 7043 9337 7049 9371
rect 7003 9249 7049 9337
rect 7261 9443 7307 9531
rect 7335 9528 7351 9580
rect 7403 9528 7423 9580
rect 7475 9528 7491 9580
rect 7261 9409 7267 9443
rect 7301 9409 7307 9443
rect 7261 9371 7307 9409
rect 7261 9337 7267 9371
rect 7301 9337 7307 9371
rect 7261 9249 7307 9337
rect 7003 9243 7307 9249
rect 7003 9209 7102 9243
rect 7136 9209 7174 9243
rect 7208 9209 7307 9243
rect 7003 9203 7307 9209
rect 7003 9141 7049 9203
rect 7261 9141 7307 9203
rect 7003 9135 7307 9141
rect 7003 9101 7102 9135
rect 7136 9101 7174 9135
rect 7208 9101 7307 9135
rect 7003 9095 7307 9101
rect 7003 9007 7049 9095
rect 7003 8973 7009 9007
rect 7043 8973 7049 9007
rect 7003 8935 7049 8973
rect 7003 8901 7009 8935
rect 7043 8901 7049 8935
rect 7003 8813 7049 8901
rect 7261 9007 7307 9095
rect 7261 8973 7267 9007
rect 7301 8973 7307 9007
rect 7261 8935 7307 8973
rect 7261 8901 7267 8935
rect 7301 8901 7307 8935
rect 7261 8813 7307 8901
rect 7519 9443 7565 9773
rect 7777 10315 7823 10645
rect 8035 10751 8081 10885
rect 8035 10717 8041 10751
rect 8075 10717 8081 10751
rect 8035 10679 8081 10717
rect 8035 10645 8041 10679
rect 8075 10645 8081 10679
rect 7851 10508 7867 10560
rect 7919 10508 7939 10560
rect 7991 10508 8007 10560
rect 7851 10400 7867 10452
rect 7919 10400 7939 10452
rect 7991 10400 8007 10452
rect 7777 10281 7783 10315
rect 7817 10281 7823 10315
rect 7777 10243 7823 10281
rect 7777 10209 7783 10243
rect 7817 10209 7823 10243
rect 7777 9879 7823 10209
rect 7777 9845 7783 9879
rect 7817 9845 7823 9879
rect 7777 9807 7823 9845
rect 7777 9773 7783 9807
rect 7817 9773 7823 9807
rect 7593 9636 7609 9688
rect 7661 9636 7681 9688
rect 7733 9636 7749 9688
rect 7593 9528 7609 9580
rect 7661 9528 7681 9580
rect 7733 9528 7749 9580
rect 7519 9409 7525 9443
rect 7559 9409 7565 9443
rect 7519 9371 7565 9409
rect 7519 9337 7525 9371
rect 7559 9337 7565 9371
rect 7519 9007 7565 9337
rect 7519 8973 7525 9007
rect 7559 8973 7565 9007
rect 7519 8935 7565 8973
rect 7519 8901 7525 8935
rect 7559 8901 7565 8935
rect 7003 8807 7307 8813
rect 7003 8773 7102 8807
rect 7136 8773 7174 8807
rect 7208 8773 7307 8807
rect 7003 8767 7307 8773
rect 7003 8705 7049 8767
rect 7261 8705 7307 8767
rect 7335 8764 7351 8816
rect 7403 8764 7423 8816
rect 7475 8764 7491 8816
rect 7003 8699 7307 8705
rect 7003 8665 7102 8699
rect 7136 8665 7174 8699
rect 7208 8665 7307 8699
rect 7003 8659 7307 8665
rect 7003 8571 7049 8659
rect 7003 8537 7009 8571
rect 7043 8537 7049 8571
rect 7003 8499 7049 8537
rect 7003 8465 7009 8499
rect 7043 8465 7049 8499
rect 7003 8377 7049 8465
rect 7261 8571 7307 8659
rect 7335 8656 7351 8708
rect 7403 8656 7423 8708
rect 7475 8656 7491 8708
rect 7261 8537 7267 8571
rect 7301 8537 7307 8571
rect 7261 8499 7307 8537
rect 7261 8465 7267 8499
rect 7301 8465 7307 8499
rect 7261 8377 7307 8465
rect 7003 8371 7307 8377
rect 7003 8337 7102 8371
rect 7136 8337 7174 8371
rect 7208 8337 7307 8371
rect 7003 8331 7307 8337
rect 7003 8269 7049 8331
rect 7261 8269 7307 8331
rect 7519 8571 7565 8901
rect 7777 9443 7823 9773
rect 8035 10315 8081 10645
rect 8293 10879 8597 10885
rect 8293 10845 8392 10879
rect 8426 10845 8464 10879
rect 8498 10845 8597 10879
rect 8293 10839 8597 10845
rect 8293 10751 8339 10839
rect 8293 10717 8299 10751
rect 8333 10717 8339 10751
rect 8293 10679 8339 10717
rect 8293 10645 8299 10679
rect 8333 10645 8339 10679
rect 8109 10508 8125 10560
rect 8177 10508 8197 10560
rect 8249 10508 8265 10560
rect 8293 10557 8339 10645
rect 8551 10751 8597 10839
rect 8551 10717 8557 10751
rect 8591 10717 8597 10751
rect 8551 10679 8597 10717
rect 8551 10645 8557 10679
rect 8591 10645 8597 10679
rect 8551 10557 8597 10645
rect 8293 10551 8597 10557
rect 8293 10517 8392 10551
rect 8426 10517 8464 10551
rect 8498 10517 8597 10551
rect 8293 10511 8597 10517
rect 8109 10400 8125 10452
rect 8177 10400 8197 10452
rect 8249 10400 8265 10452
rect 8293 10449 8339 10511
rect 8551 10449 8597 10511
rect 9916 10829 10178 10877
rect 9916 10777 10024 10829
rect 10076 10777 10178 10829
rect 9916 10456 10178 10777
rect 8293 10443 8597 10449
rect 8293 10409 8392 10443
rect 8426 10409 8464 10443
rect 8498 10409 8597 10443
rect 8293 10403 8597 10409
rect 8035 10281 8041 10315
rect 8075 10281 8081 10315
rect 8035 10243 8081 10281
rect 8035 10209 8041 10243
rect 8075 10209 8081 10243
rect 8035 9879 8081 10209
rect 8035 9845 8041 9879
rect 8075 9845 8081 9879
rect 8035 9807 8081 9845
rect 8035 9773 8041 9807
rect 8075 9773 8081 9807
rect 7851 9636 7867 9688
rect 7919 9636 7939 9688
rect 7991 9636 8007 9688
rect 7851 9528 7867 9580
rect 7919 9528 7939 9580
rect 7991 9528 8007 9580
rect 7777 9409 7783 9443
rect 7817 9409 7823 9443
rect 7777 9371 7823 9409
rect 7777 9337 7783 9371
rect 7817 9337 7823 9371
rect 7777 9007 7823 9337
rect 7777 8973 7783 9007
rect 7817 8973 7823 9007
rect 7777 8935 7823 8973
rect 7777 8901 7783 8935
rect 7817 8901 7823 8935
rect 7593 8764 7609 8816
rect 7661 8764 7681 8816
rect 7733 8764 7749 8816
rect 7593 8656 7609 8708
rect 7661 8656 7681 8708
rect 7733 8656 7749 8708
rect 7519 8537 7525 8571
rect 7559 8537 7565 8571
rect 7519 8499 7565 8537
rect 7519 8465 7525 8499
rect 7559 8465 7565 8499
rect 7003 8263 7307 8269
rect 7003 8229 7102 8263
rect 7136 8229 7174 8263
rect 7208 8229 7307 8263
rect 7003 8223 7307 8229
rect 7003 8135 7049 8223
rect 7003 8101 7009 8135
rect 7043 8101 7049 8135
rect 7003 8063 7049 8101
rect 7003 8029 7009 8063
rect 7043 8029 7049 8063
rect 670 7979 1186 7982
rect -1956 7903 -1910 7979
rect -1956 7869 -1950 7903
rect -1916 7869 -1910 7903
rect -1956 7831 -1910 7869
rect -1956 7797 -1950 7831
rect -1916 7797 -1910 7831
rect -1956 7718 -1910 7797
rect -2214 7712 -1910 7718
rect -2214 7678 -2115 7712
rect -2081 7678 -2043 7712
rect -2009 7678 -1910 7712
rect -2214 7672 -1910 7678
rect -2214 7610 -2168 7672
rect -1956 7613 -1910 7672
rect -1701 7903 -1649 7979
rect -1701 7869 -1692 7903
rect -1658 7869 -1649 7903
rect -1701 7831 -1649 7869
rect -1701 7797 -1692 7831
rect -1658 7797 -1649 7831
rect -1701 7613 -1649 7797
rect -1440 7903 -1394 7979
rect -1440 7869 -1434 7903
rect -1400 7869 -1394 7903
rect -1440 7831 -1394 7869
rect -1440 7797 -1434 7831
rect -1400 7797 -1394 7831
rect -1440 7750 -1394 7797
rect -1185 7903 -1133 7979
rect -1185 7869 -1176 7903
rect -1142 7869 -1133 7903
rect -1185 7831 -1133 7869
rect -1185 7797 -1176 7831
rect -1142 7797 -1133 7831
rect -1185 7750 -1133 7797
rect -924 7903 -878 7950
rect -924 7869 -918 7903
rect -884 7869 -878 7903
rect -924 7831 -878 7869
rect -924 7797 -918 7831
rect -884 7797 -878 7831
rect -1956 7610 -1440 7613
rect -2214 7604 -1440 7610
rect -2214 7570 -2115 7604
rect -2081 7570 -2043 7604
rect -2009 7570 -1857 7604
rect -1823 7570 -1785 7604
rect -1751 7570 -1599 7604
rect -1565 7570 -1527 7604
rect -1493 7570 -1440 7604
rect -2214 7564 -1440 7570
rect -2214 7485 -2168 7564
rect -2214 7451 -2208 7485
rect -2174 7451 -2168 7485
rect -2214 7413 -2168 7451
rect -2214 7379 -2208 7413
rect -2174 7379 -2168 7413
rect -2214 7300 -2168 7379
rect -1956 7561 -1440 7564
rect -1366 7561 -1350 7613
rect -1298 7561 -1278 7613
rect -1226 7561 -1192 7613
rect -1126 7561 -1092 7613
rect -1040 7561 -1020 7613
rect -968 7561 -952 7613
rect -1956 7485 -1910 7561
rect -1956 7451 -1950 7485
rect -1916 7451 -1910 7485
rect -1956 7413 -1910 7451
rect -1956 7379 -1950 7413
rect -1916 7379 -1910 7413
rect -1956 7300 -1910 7379
rect -1701 7485 -1649 7561
rect -1701 7451 -1692 7485
rect -1658 7451 -1649 7485
rect -1701 7413 -1649 7451
rect -1701 7379 -1692 7413
rect -1658 7379 -1649 7413
rect -1701 7332 -1649 7379
rect -1440 7485 -1394 7532
rect -1440 7451 -1434 7485
rect -1400 7451 -1394 7485
rect -1440 7413 -1394 7451
rect -1440 7379 -1434 7413
rect -1400 7379 -1394 7413
rect -2214 7294 -1910 7300
rect -2214 7260 -2115 7294
rect -2081 7260 -2043 7294
rect -2009 7260 -1910 7294
rect -2214 7254 -1910 7260
rect -1440 7272 -1394 7379
rect -1185 7494 -1133 7532
rect -1185 7422 -1133 7442
rect -1185 7332 -1133 7370
rect -924 7485 -878 7797
rect -669 7912 -617 7950
rect -669 7840 -617 7860
rect -669 7750 -617 7788
rect -408 7903 -362 7950
rect -408 7869 -402 7903
rect -368 7869 -362 7903
rect -408 7831 -362 7869
rect -408 7797 -402 7831
rect -368 7797 -362 7831
rect -924 7451 -918 7485
rect -884 7451 -878 7485
rect -924 7413 -878 7451
rect -924 7379 -918 7413
rect -884 7379 -878 7413
rect -924 7272 -878 7379
rect -669 7494 -617 7532
rect -669 7422 -617 7442
rect -669 7332 -617 7370
rect -408 7485 -362 7797
rect -153 7912 -101 7950
rect -153 7840 -101 7860
rect -153 7750 -101 7788
rect 108 7903 154 7950
rect 108 7869 114 7903
rect 148 7869 154 7903
rect 108 7831 154 7869
rect 108 7797 114 7831
rect 148 7797 154 7831
rect -334 7561 -318 7613
rect -266 7561 -246 7613
rect -194 7561 -160 7613
rect -94 7561 -60 7613
rect -8 7561 12 7613
rect 64 7561 80 7613
rect -408 7451 -402 7485
rect -368 7451 -362 7485
rect -408 7413 -362 7451
rect -408 7379 -402 7413
rect -368 7379 -362 7413
rect -2214 7192 -2168 7254
rect -1440 7226 -878 7272
rect -850 7251 -834 7303
rect -782 7251 -762 7303
rect -710 7251 -676 7303
rect -610 7251 -576 7303
rect -524 7251 -504 7303
rect -452 7251 -436 7303
rect -408 7274 -362 7379
rect -153 7494 -101 7532
rect -153 7422 -101 7442
rect -153 7332 -101 7370
rect 108 7485 154 7797
rect 363 7912 415 7950
rect 363 7840 415 7860
rect 363 7750 415 7788
rect 624 7903 670 7950
rect 624 7869 630 7903
rect 664 7869 670 7903
rect 624 7831 670 7869
rect 624 7797 630 7831
rect 664 7797 670 7831
rect 108 7451 114 7485
rect 148 7451 154 7485
rect 108 7413 154 7451
rect 108 7379 114 7413
rect 148 7379 154 7413
rect 108 7274 154 7379
rect 363 7494 415 7532
rect 363 7422 415 7442
rect 363 7332 415 7370
rect 624 7485 670 7797
rect 879 7903 931 7979
rect 879 7869 888 7903
rect 922 7869 931 7903
rect 879 7831 931 7869
rect 879 7797 888 7831
rect 922 7797 931 7831
rect 879 7750 931 7797
rect 1140 7903 1186 7979
rect 1140 7869 1146 7903
rect 1180 7869 1186 7903
rect 1140 7831 1186 7869
rect 1140 7797 1146 7831
rect 1180 7797 1186 7831
rect 1140 7750 1186 7797
rect 1398 7903 1444 7982
rect 3197 7930 3211 7982
rect 3263 7930 5187 7982
rect 7003 7941 7049 8029
rect 7261 8135 7307 8223
rect 7335 8220 7351 8272
rect 7403 8220 7423 8272
rect 7475 8220 7491 8272
rect 7261 8101 7267 8135
rect 7301 8101 7307 8135
rect 7261 8063 7307 8101
rect 7261 8029 7267 8063
rect 7301 8029 7307 8063
rect 7261 7941 7307 8029
rect 7003 7935 7307 7941
rect 1398 7869 1404 7903
rect 1438 7869 1444 7903
rect 7003 7901 7102 7935
rect 7136 7901 7174 7935
rect 7208 7901 7307 7935
rect 7003 7895 7307 7901
rect 7519 8135 7565 8465
rect 7777 8571 7823 8901
rect 8035 9443 8081 9773
rect 8293 10315 8339 10403
rect 8293 10281 8299 10315
rect 8333 10281 8339 10315
rect 8293 10243 8339 10281
rect 8293 10209 8299 10243
rect 8333 10209 8339 10243
rect 8293 10121 8339 10209
rect 8551 10315 8597 10403
rect 8551 10281 8557 10315
rect 8591 10281 8597 10315
rect 8551 10243 8597 10281
rect 8551 10209 8557 10243
rect 8591 10209 8597 10243
rect 8551 10121 8597 10209
rect 8293 10115 8597 10121
rect 8293 10081 8392 10115
rect 8426 10081 8464 10115
rect 8498 10081 8597 10115
rect 8293 10075 8597 10081
rect 8293 10013 8339 10075
rect 8551 10013 8597 10075
rect 8293 10007 8597 10013
rect 8293 9973 8392 10007
rect 8426 9973 8464 10007
rect 8498 9973 8597 10007
rect 8293 9967 8597 9973
rect 8293 9879 8339 9967
rect 8293 9845 8299 9879
rect 8333 9845 8339 9879
rect 8293 9807 8339 9845
rect 8293 9773 8299 9807
rect 8333 9773 8339 9807
rect 8109 9636 8125 9688
rect 8177 9636 8197 9688
rect 8249 9636 8265 9688
rect 8293 9685 8339 9773
rect 8551 9879 8597 9967
rect 8551 9845 8557 9879
rect 8591 9845 8597 9879
rect 8551 9807 8597 9845
rect 8551 9773 8557 9807
rect 8591 9773 8597 9807
rect 8551 9685 8597 9773
rect 8293 9679 8597 9685
rect 8293 9645 8392 9679
rect 8426 9645 8464 9679
rect 8498 9645 8597 9679
rect 8293 9639 8597 9645
rect 8109 9528 8125 9580
rect 8177 9528 8197 9580
rect 8249 9528 8265 9580
rect 8293 9577 8339 9639
rect 8551 9577 8597 9639
rect 8293 9571 8597 9577
rect 8293 9537 8392 9571
rect 8426 9537 8464 9571
rect 8498 9537 8597 9571
rect 8293 9531 8597 9537
rect 8035 9409 8041 9443
rect 8075 9409 8081 9443
rect 8035 9371 8081 9409
rect 8035 9337 8041 9371
rect 8075 9337 8081 9371
rect 8035 9007 8081 9337
rect 8035 8973 8041 9007
rect 8075 8973 8081 9007
rect 8035 8935 8081 8973
rect 8035 8901 8041 8935
rect 8075 8901 8081 8935
rect 7851 8764 7867 8816
rect 7919 8764 7939 8816
rect 7991 8764 8007 8816
rect 7851 8656 7867 8708
rect 7919 8656 7939 8708
rect 7991 8656 8007 8708
rect 7777 8537 7783 8571
rect 7817 8537 7823 8571
rect 7777 8499 7823 8537
rect 7777 8465 7783 8499
rect 7817 8465 7823 8499
rect 7593 8220 7609 8272
rect 7661 8220 7681 8272
rect 7733 8220 7749 8272
rect 7519 8101 7525 8135
rect 7559 8101 7565 8135
rect 7519 8063 7565 8101
rect 7519 8029 7525 8063
rect 7559 8029 7565 8063
rect 1398 7831 1444 7869
rect 1398 7797 1404 7831
rect 1438 7797 1444 7831
rect 1398 7718 1444 7797
rect 1186 7712 1444 7718
rect 1186 7678 1239 7712
rect 1273 7678 1311 7712
rect 1345 7678 1444 7712
rect 1186 7672 1444 7678
rect 698 7561 714 7613
rect 766 7561 786 7613
rect 838 7561 872 7613
rect 938 7561 972 7613
rect 1024 7561 1044 7613
rect 1096 7561 1112 7613
rect 1398 7610 1444 7672
rect 624 7451 630 7485
rect 664 7451 670 7485
rect 624 7413 670 7451
rect 624 7379 630 7413
rect 664 7379 670 7413
rect -2214 7186 -1984 7192
rect -2214 7152 -2115 7186
rect -2081 7152 -2043 7186
rect -2009 7152 -1984 7186
rect -2214 7146 -1984 7152
rect -2214 7067 -2168 7146
rect -2214 7033 -2208 7067
rect -2174 7033 -2168 7067
rect -2214 6995 -2168 7033
rect -2214 6961 -2208 6995
rect -2174 6961 -2168 6995
rect -2214 6882 -2168 6961
rect -1956 7067 -1910 7192
rect -1882 7143 -1866 7195
rect -1814 7143 -1794 7195
rect -1742 7143 -1708 7195
rect -1642 7143 -1608 7195
rect -1556 7143 -1536 7195
rect -1484 7143 -1468 7195
rect -1956 7033 -1950 7067
rect -1916 7033 -1910 7067
rect -1956 6995 -1910 7033
rect -1956 6961 -1950 6995
rect -1916 6961 -1910 6995
rect -2214 6876 -1984 6882
rect -2214 6842 -2115 6876
rect -2081 6842 -2043 6876
rect -2009 6842 -1984 6876
rect -2214 6836 -1984 6842
rect -2214 6774 -2168 6836
rect -1956 6816 -1910 6961
rect -1701 7076 -1649 7114
rect -1701 7004 -1649 7024
rect -1701 6914 -1649 6952
rect -1440 7067 -1394 7226
rect -1440 7033 -1434 7067
rect -1400 7033 -1394 7067
rect -1440 6995 -1394 7033
rect -1440 6961 -1434 6995
rect -1400 6961 -1394 6995
rect -1440 6816 -1394 6961
rect -1185 7076 -1133 7114
rect -1185 7004 -1133 7024
rect -1185 6914 -1133 6952
rect -924 7067 -878 7226
rect -408 7228 154 7274
rect 182 7251 198 7303
rect 250 7251 270 7303
rect 322 7251 356 7303
rect 422 7251 456 7303
rect 508 7251 528 7303
rect 580 7251 596 7303
rect 624 7279 670 7379
rect 879 7494 931 7532
rect 879 7422 931 7442
rect 879 7332 931 7370
rect 1140 7485 1186 7610
rect 1214 7604 1444 7610
rect 1214 7570 1239 7604
rect 1273 7570 1311 7604
rect 1345 7570 1444 7604
rect 1214 7564 1444 7570
rect 7519 7567 7565 8029
rect 7777 8135 7823 8465
rect 8035 8571 8081 8901
rect 8293 9443 8339 9531
rect 8293 9409 8299 9443
rect 8333 9409 8339 9443
rect 8293 9371 8339 9409
rect 8293 9337 8299 9371
rect 8333 9337 8339 9371
rect 8293 9249 8339 9337
rect 8551 9443 8597 9531
rect 8551 9409 8557 9443
rect 8591 9409 8597 9443
rect 8551 9371 8597 9409
rect 8551 9337 8557 9371
rect 8591 9337 8597 9371
rect 8551 9249 8597 9337
rect 8293 9243 8597 9249
rect 8293 9209 8392 9243
rect 8426 9209 8464 9243
rect 8498 9209 8597 9243
rect 8293 9203 8597 9209
rect 8293 9141 8339 9203
rect 8551 9141 8597 9203
rect 8293 9135 8597 9141
rect 8293 9101 8392 9135
rect 8426 9101 8464 9135
rect 8498 9101 8597 9135
rect 8293 9095 8597 9101
rect 8293 9007 8339 9095
rect 8293 8973 8299 9007
rect 8333 8973 8339 9007
rect 8293 8935 8339 8973
rect 8293 8901 8299 8935
rect 8333 8901 8339 8935
rect 8109 8764 8125 8816
rect 8177 8764 8197 8816
rect 8249 8764 8265 8816
rect 8293 8813 8339 8901
rect 8551 9007 8597 9095
rect 8551 8973 8557 9007
rect 8591 8973 8597 9007
rect 8551 8935 8597 8973
rect 8551 8901 8557 8935
rect 8591 8901 8597 8935
rect 8551 8813 8597 8901
rect 8293 8807 8597 8813
rect 8293 8773 8392 8807
rect 8426 8773 8464 8807
rect 8498 8773 8597 8807
rect 8293 8767 8597 8773
rect 8109 8656 8125 8708
rect 8177 8656 8197 8708
rect 8249 8656 8265 8708
rect 8293 8705 8339 8767
rect 8551 8705 8597 8767
rect 8293 8699 8597 8705
rect 8293 8665 8392 8699
rect 8426 8665 8464 8699
rect 8498 8665 8597 8699
rect 8293 8659 8597 8665
rect 8035 8537 8041 8571
rect 8075 8537 8081 8571
rect 8035 8499 8081 8537
rect 8035 8465 8041 8499
rect 8075 8465 8081 8499
rect 7851 8220 7867 8272
rect 7919 8220 7939 8272
rect 7991 8220 8007 8272
rect 7777 8101 7783 8135
rect 7817 8101 7823 8135
rect 7777 8063 7823 8101
rect 7777 8029 7783 8063
rect 7817 8029 7823 8063
rect 7777 7895 7823 8029
rect 8035 8135 8081 8465
rect 8293 8571 8339 8659
rect 8293 8537 8299 8571
rect 8333 8537 8339 8571
rect 8293 8499 8339 8537
rect 8293 8465 8299 8499
rect 8333 8465 8339 8499
rect 8293 8377 8339 8465
rect 8551 8571 8597 8659
rect 8551 8537 8557 8571
rect 8591 8537 8597 8571
rect 8551 8499 8597 8537
rect 8551 8465 8557 8499
rect 8591 8465 8597 8499
rect 8551 8377 8597 8465
rect 8293 8371 8597 8377
rect 8293 8337 8392 8371
rect 8426 8337 8464 8371
rect 8498 8337 8597 8371
rect 8293 8331 8597 8337
rect 8109 8220 8125 8272
rect 8177 8220 8197 8272
rect 8249 8220 8265 8272
rect 8293 8269 8339 8331
rect 8551 8269 8597 8331
rect 8293 8263 8597 8269
rect 8293 8229 8392 8263
rect 8426 8229 8464 8263
rect 8498 8229 8597 8263
rect 8293 8223 8597 8229
rect 8035 8101 8041 8135
rect 8075 8101 8081 8135
rect 8035 8063 8081 8101
rect 8035 8029 8041 8063
rect 8075 8029 8081 8063
rect 8035 7567 8081 8029
rect 8293 8135 8339 8223
rect 8293 8101 8299 8135
rect 8333 8101 8339 8135
rect 8293 8063 8339 8101
rect 8293 8029 8299 8063
rect 8333 8029 8339 8063
rect 8293 7941 8339 8029
rect 8551 8135 8597 8223
rect 8551 8101 8557 8135
rect 8591 8101 8597 8135
rect 8551 8063 8597 8101
rect 8551 8029 8557 8063
rect 8591 8029 8597 8063
rect 8551 7941 8597 8029
rect 8293 7935 8597 7941
rect 8293 7901 8392 7935
rect 8426 7901 8464 7935
rect 8498 7901 8597 7935
rect 8293 7895 8597 7901
rect 9583 8511 12333 8557
rect 9583 7567 9629 8511
rect 9916 8146 10178 8278
rect 9916 8064 10861 8146
rect 9916 8004 11163 8064
rect 9916 7986 10861 8004
rect 9916 7857 10178 7986
rect 1140 7451 1146 7485
rect 1180 7451 1186 7485
rect 1140 7413 1186 7451
rect 1140 7379 1146 7413
rect 1180 7379 1186 7413
rect 1140 7279 1186 7379
rect 1398 7485 1444 7564
rect 7003 7521 9629 7567
rect 9893 7605 10333 7658
rect 1398 7451 1404 7485
rect 1438 7451 1444 7485
rect 1398 7413 1444 7451
rect 1398 7379 1404 7413
rect 1438 7379 1444 7413
rect 1398 7300 1444 7379
rect -850 7143 -834 7195
rect -782 7143 -762 7195
rect -710 7143 -676 7195
rect -610 7143 -576 7195
rect -524 7143 -504 7195
rect -452 7143 -436 7195
rect -924 7033 -918 7067
rect -884 7033 -878 7067
rect -924 6995 -878 7033
rect -924 6961 -918 6995
rect -884 6961 -878 6995
rect -1366 6833 -1350 6885
rect -1298 6833 -1278 6885
rect -1226 6833 -1192 6885
rect -1126 6833 -1092 6885
rect -1040 6833 -1020 6885
rect -968 6833 -952 6885
rect -2214 6768 -1984 6774
rect -2214 6734 -2115 6768
rect -2081 6734 -2043 6768
rect -2009 6734 -1984 6768
rect -2214 6728 -1984 6734
rect -1956 6770 -1394 6816
rect -924 6805 -878 6961
rect -669 7076 -617 7114
rect -669 7004 -617 7024
rect -669 6914 -617 6952
rect -408 7067 -362 7228
rect -408 7033 -402 7067
rect -368 7033 -362 7067
rect -408 6995 -362 7033
rect -408 6961 -402 6995
rect -368 6961 -362 6995
rect -408 6805 -362 6961
rect -153 7076 -101 7114
rect -153 7004 -101 7024
rect -153 6914 -101 6952
rect 108 7067 154 7228
rect 624 7233 1186 7279
rect 1214 7294 1444 7300
rect 1214 7260 1239 7294
rect 1273 7260 1311 7294
rect 1345 7260 1444 7294
rect 1214 7254 1444 7260
rect 182 7143 198 7195
rect 250 7143 270 7195
rect 322 7143 356 7195
rect 422 7143 456 7195
rect 508 7143 528 7195
rect 580 7143 596 7195
rect 108 7033 114 7067
rect 148 7033 154 7067
rect 108 6995 154 7033
rect 108 6961 114 6995
rect 148 6961 154 6995
rect -334 6833 -318 6885
rect -266 6833 -246 6885
rect -194 6833 -160 6885
rect -94 6833 -60 6885
rect -8 6833 12 6885
rect 64 6833 80 6885
rect -2214 6649 -2168 6728
rect -2214 6615 -2208 6649
rect -2174 6615 -2168 6649
rect -2214 6577 -2168 6615
rect -2214 6543 -2208 6577
rect -2174 6543 -2168 6577
rect -2214 6464 -2168 6543
rect -1956 6649 -1910 6770
rect -1956 6615 -1950 6649
rect -1916 6615 -1910 6649
rect -1956 6577 -1910 6615
rect -1956 6543 -1950 6577
rect -1916 6543 -1910 6577
rect -2214 6458 -1984 6464
rect -2214 6424 -2115 6458
rect -2081 6424 -2043 6458
rect -2009 6424 -1984 6458
rect -2214 6418 -1984 6424
rect -2214 6356 -2168 6418
rect -2214 6350 -1984 6356
rect -2214 6316 -2115 6350
rect -2081 6316 -2043 6350
rect -2009 6316 -1984 6350
rect -2214 6310 -1984 6316
rect -2214 6231 -2168 6310
rect -2214 6197 -2208 6231
rect -2174 6197 -2168 6231
rect -2214 6159 -2168 6197
rect -2214 6125 -2208 6159
rect -2174 6125 -2168 6159
rect -2214 6046 -2168 6125
rect -1956 6231 -1910 6543
rect -1701 6658 -1649 6696
rect -1701 6586 -1649 6606
rect -1701 6496 -1649 6534
rect -1440 6649 -1394 6770
rect -1366 6725 -1350 6777
rect -1298 6725 -1278 6777
rect -1226 6725 -1192 6777
rect -1126 6725 -1092 6777
rect -1040 6725 -1020 6777
rect -968 6725 -952 6777
rect -924 6759 -362 6805
rect 108 6800 154 6961
rect 363 7076 415 7114
rect 363 7004 415 7024
rect 363 6914 415 6952
rect 624 7067 670 7233
rect 624 7033 630 7067
rect 664 7033 670 7067
rect 624 6995 670 7033
rect 624 6961 630 6995
rect 664 6961 670 6995
rect 624 6800 670 6961
rect 879 7076 931 7114
rect 879 7004 931 7024
rect 879 6914 931 6952
rect 1140 7067 1186 7233
rect 1398 7192 1444 7254
rect 1214 7186 1444 7192
rect 1214 7152 1239 7186
rect 1273 7152 1311 7186
rect 1345 7152 1444 7186
rect 1214 7146 1444 7152
rect 1140 7033 1146 7067
rect 1180 7033 1186 7067
rect 1140 6995 1186 7033
rect 1140 6961 1146 6995
rect 1180 6961 1186 6995
rect 698 6833 714 6885
rect 766 6833 786 6885
rect 838 6833 872 6885
rect 938 6833 972 6885
rect 1024 6833 1044 6885
rect 1096 6833 1112 6885
rect -1440 6615 -1434 6649
rect -1400 6615 -1394 6649
rect -1440 6577 -1394 6615
rect -1440 6543 -1434 6577
rect -1400 6543 -1394 6577
rect -1882 6415 -1866 6467
rect -1814 6415 -1794 6467
rect -1742 6415 -1708 6467
rect -1642 6415 -1608 6467
rect -1556 6415 -1536 6467
rect -1484 6415 -1468 6467
rect -1882 6307 -1866 6359
rect -1814 6307 -1794 6359
rect -1742 6307 -1708 6359
rect -1642 6307 -1608 6359
rect -1556 6307 -1536 6359
rect -1484 6307 -1468 6359
rect -1956 6197 -1950 6231
rect -1916 6197 -1910 6231
rect -1956 6159 -1910 6197
rect -1956 6125 -1950 6159
rect -1916 6125 -1910 6159
rect -2214 6040 -1984 6046
rect -2214 6006 -2115 6040
rect -2081 6006 -2043 6040
rect -2009 6006 -1984 6040
rect -2214 6000 -1984 6006
rect -2214 5938 -2168 6000
rect -2214 5932 -1984 5938
rect -2214 5898 -2115 5932
rect -2081 5898 -2043 5932
rect -2009 5898 -1984 5932
rect -2214 5892 -1984 5898
rect -2214 5813 -2168 5892
rect -2214 5779 -2208 5813
rect -2174 5779 -2168 5813
rect -2214 5741 -2168 5779
rect -2214 5707 -2208 5741
rect -2174 5707 -2168 5741
rect -2214 5628 -2168 5707
rect -1956 5813 -1910 6125
rect -1701 6240 -1649 6278
rect -1701 6168 -1649 6188
rect -1701 6078 -1649 6116
rect -1440 6231 -1394 6543
rect -1185 6658 -1133 6696
rect -1185 6586 -1133 6606
rect -1185 6496 -1133 6534
rect -924 6649 -878 6759
rect -924 6615 -918 6649
rect -884 6615 -878 6649
rect -924 6577 -878 6615
rect -924 6543 -918 6577
rect -884 6543 -878 6577
rect -1440 6197 -1434 6231
rect -1400 6197 -1394 6231
rect -1440 6159 -1394 6197
rect -1440 6125 -1434 6159
rect -1400 6125 -1394 6159
rect -1956 5779 -1950 5813
rect -1916 5779 -1910 5813
rect -1956 5741 -1910 5779
rect -1956 5707 -1950 5741
rect -1916 5707 -1910 5741
rect -2214 5622 -1984 5628
rect -2214 5588 -2115 5622
rect -2081 5588 -2043 5622
rect -2009 5588 -1984 5622
rect -2214 5582 -1984 5588
rect -2214 5520 -2168 5582
rect -2214 5514 -1984 5520
rect -2214 5480 -2115 5514
rect -2081 5480 -2043 5514
rect -2009 5480 -1984 5514
rect -2214 5474 -1984 5480
rect -2214 5395 -2168 5474
rect -2214 5361 -2208 5395
rect -2174 5361 -2168 5395
rect -2214 5323 -2168 5361
rect -2214 5289 -2208 5323
rect -2174 5289 -2168 5323
rect -2214 5210 -2168 5289
rect -1956 5395 -1910 5707
rect -1701 5822 -1649 5860
rect -1701 5750 -1649 5770
rect -1701 5660 -1649 5698
rect -1440 5813 -1394 6125
rect -1185 6240 -1133 6278
rect -1185 6168 -1133 6188
rect -1185 6078 -1133 6116
rect -924 6231 -878 6543
rect -669 6658 -617 6696
rect -669 6586 -617 6606
rect -669 6496 -617 6534
rect -408 6649 -362 6759
rect -334 6725 -318 6777
rect -266 6725 -246 6777
rect -194 6725 -160 6777
rect -94 6725 -60 6777
rect -8 6725 12 6777
rect 64 6725 80 6777
rect 108 6754 670 6800
rect -408 6615 -402 6649
rect -368 6615 -362 6649
rect -408 6577 -362 6615
rect -408 6543 -402 6577
rect -368 6543 -362 6577
rect -850 6415 -834 6467
rect -782 6415 -762 6467
rect -710 6415 -676 6467
rect -610 6415 -576 6467
rect -524 6415 -504 6467
rect -452 6415 -436 6467
rect -850 6307 -834 6359
rect -782 6307 -762 6359
rect -710 6307 -676 6359
rect -610 6307 -576 6359
rect -524 6307 -504 6359
rect -452 6307 -436 6359
rect -924 6197 -918 6231
rect -884 6197 -878 6231
rect -924 6159 -878 6197
rect -924 6125 -918 6159
rect -884 6125 -878 6159
rect -1366 5997 -1350 6049
rect -1298 5997 -1278 6049
rect -1226 5997 -1192 6049
rect -1126 5997 -1092 6049
rect -1040 5997 -1020 6049
rect -968 5997 -952 6049
rect -1366 5889 -1350 5941
rect -1298 5889 -1278 5941
rect -1226 5889 -1192 5941
rect -1126 5889 -1092 5941
rect -1040 5889 -1020 5941
rect -968 5889 -952 5941
rect -1440 5779 -1434 5813
rect -1400 5779 -1394 5813
rect -1440 5741 -1394 5779
rect -1440 5707 -1434 5741
rect -1400 5707 -1394 5741
rect -1882 5579 -1866 5631
rect -1814 5579 -1794 5631
rect -1742 5579 -1708 5631
rect -1642 5579 -1608 5631
rect -1556 5579 -1536 5631
rect -1484 5579 -1468 5631
rect -1882 5471 -1866 5523
rect -1814 5471 -1794 5523
rect -1742 5471 -1708 5523
rect -1642 5471 -1608 5523
rect -1556 5471 -1536 5523
rect -1484 5471 -1468 5523
rect -1956 5361 -1950 5395
rect -1916 5361 -1910 5395
rect -1956 5323 -1910 5361
rect -1956 5289 -1950 5323
rect -1916 5289 -1910 5323
rect -2214 5204 -1984 5210
rect -2214 5170 -2115 5204
rect -2081 5170 -2043 5204
rect -2009 5170 -1984 5204
rect -2214 5164 -1984 5170
rect -2214 5102 -2168 5164
rect -2214 5096 -1984 5102
rect -2214 5062 -2115 5096
rect -2081 5062 -2043 5096
rect -2009 5062 -1984 5096
rect -2214 5056 -1984 5062
rect -2214 4977 -2168 5056
rect -2214 4943 -2208 4977
rect -2174 4943 -2168 4977
rect -2214 4905 -2168 4943
rect -2214 4871 -2208 4905
rect -2174 4871 -2168 4905
rect -2214 4792 -2168 4871
rect -1956 4977 -1910 5289
rect -1701 5404 -1649 5442
rect -1701 5332 -1649 5352
rect -1701 5242 -1649 5280
rect -1440 5395 -1394 5707
rect -1185 5822 -1133 5860
rect -1185 5750 -1133 5770
rect -1185 5660 -1133 5698
rect -924 5813 -878 6125
rect -669 6240 -617 6278
rect -669 6168 -617 6188
rect -669 6078 -617 6116
rect -408 6231 -362 6543
rect -153 6658 -101 6696
rect -153 6586 -101 6606
rect -153 6496 -101 6534
rect 108 6649 154 6754
rect 108 6615 114 6649
rect 148 6615 154 6649
rect 108 6577 154 6615
rect 108 6543 114 6577
rect 148 6543 154 6577
rect -408 6197 -402 6231
rect -368 6197 -362 6231
rect -408 6159 -362 6197
rect -408 6125 -402 6159
rect -368 6125 -362 6159
rect -924 5779 -918 5813
rect -884 5779 -878 5813
rect -924 5741 -878 5779
rect -924 5707 -918 5741
rect -884 5707 -878 5741
rect -1440 5361 -1434 5395
rect -1400 5361 -1394 5395
rect -1440 5323 -1394 5361
rect -1440 5289 -1434 5323
rect -1400 5289 -1394 5323
rect -1956 4943 -1950 4977
rect -1916 4943 -1910 4977
rect -1956 4905 -1910 4943
rect -1956 4871 -1950 4905
rect -1916 4871 -1910 4905
rect -2214 4786 -1984 4792
rect -2214 4752 -2115 4786
rect -2081 4752 -2043 4786
rect -2009 4752 -1984 4786
rect -2214 4746 -1984 4752
rect -2214 4684 -2168 4746
rect -2214 4678 -1984 4684
rect -2214 4644 -2115 4678
rect -2081 4644 -2043 4678
rect -2009 4644 -1984 4678
rect -2214 4638 -1984 4644
rect -2214 4559 -2168 4638
rect -2214 4525 -2208 4559
rect -2174 4525 -2168 4559
rect -2214 4487 -2168 4525
rect -2214 4453 -2208 4487
rect -2174 4453 -2168 4487
rect -2214 4374 -2168 4453
rect -1956 4559 -1910 4871
rect -1701 4986 -1649 5024
rect -1701 4914 -1649 4934
rect -1701 4824 -1649 4862
rect -1440 4977 -1394 5289
rect -1185 5404 -1133 5442
rect -1185 5332 -1133 5352
rect -1185 5242 -1133 5280
rect -924 5395 -878 5707
rect -669 5822 -617 5860
rect -669 5750 -617 5770
rect -669 5660 -617 5698
rect -408 5813 -362 6125
rect -153 6240 -101 6278
rect -153 6168 -101 6188
rect -153 6078 -101 6116
rect 108 6231 154 6543
rect 363 6658 415 6696
rect 363 6586 415 6606
rect 363 6496 415 6534
rect 624 6649 670 6754
rect 698 6725 714 6777
rect 766 6725 786 6777
rect 838 6725 872 6777
rect 938 6725 972 6777
rect 1024 6725 1044 6777
rect 1096 6725 1112 6777
rect 624 6615 630 6649
rect 664 6615 670 6649
rect 624 6577 670 6615
rect 624 6543 630 6577
rect 664 6543 670 6577
rect 182 6415 198 6467
rect 250 6415 270 6467
rect 322 6415 356 6467
rect 422 6415 456 6467
rect 508 6415 528 6467
rect 580 6415 596 6467
rect 182 6307 198 6359
rect 250 6307 270 6359
rect 322 6307 356 6359
rect 422 6307 456 6359
rect 508 6307 528 6359
rect 580 6307 596 6359
rect 108 6197 114 6231
rect 148 6197 154 6231
rect 108 6159 154 6197
rect 108 6125 114 6159
rect 148 6125 154 6159
rect -334 5997 -318 6049
rect -266 5997 -246 6049
rect -194 5997 -160 6049
rect -94 5997 -60 6049
rect -8 5997 12 6049
rect 64 5997 80 6049
rect -334 5889 -318 5941
rect -266 5889 -246 5941
rect -194 5889 -160 5941
rect -94 5889 -60 5941
rect -8 5889 12 5941
rect 64 5889 80 5941
rect -408 5779 -402 5813
rect -368 5779 -362 5813
rect -408 5741 -362 5779
rect -408 5707 -402 5741
rect -368 5707 -362 5741
rect -850 5579 -834 5631
rect -782 5579 -762 5631
rect -710 5579 -676 5631
rect -610 5579 -576 5631
rect -524 5579 -504 5631
rect -452 5579 -436 5631
rect -850 5471 -834 5523
rect -782 5471 -762 5523
rect -710 5471 -676 5523
rect -610 5471 -576 5523
rect -524 5471 -504 5523
rect -452 5471 -436 5523
rect -924 5361 -918 5395
rect -884 5361 -878 5395
rect -924 5323 -878 5361
rect -924 5289 -918 5323
rect -884 5289 -878 5323
rect -1366 5161 -1350 5213
rect -1298 5161 -1278 5213
rect -1226 5161 -1192 5213
rect -1126 5161 -1092 5213
rect -1040 5161 -1020 5213
rect -968 5161 -952 5213
rect -1366 5053 -1350 5105
rect -1298 5053 -1278 5105
rect -1226 5053 -1192 5105
rect -1126 5053 -1092 5105
rect -1040 5053 -1020 5105
rect -968 5053 -952 5105
rect -1440 4943 -1434 4977
rect -1400 4943 -1394 4977
rect -1440 4905 -1394 4943
rect -1440 4871 -1434 4905
rect -1400 4871 -1394 4905
rect -1882 4743 -1866 4795
rect -1814 4743 -1794 4795
rect -1742 4743 -1708 4795
rect -1642 4743 -1608 4795
rect -1556 4743 -1536 4795
rect -1484 4743 -1468 4795
rect -1882 4635 -1866 4687
rect -1814 4635 -1794 4687
rect -1742 4635 -1708 4687
rect -1642 4635 -1608 4687
rect -1556 4635 -1536 4687
rect -1484 4635 -1468 4687
rect -1956 4525 -1950 4559
rect -1916 4525 -1910 4559
rect -1956 4487 -1910 4525
rect -1956 4453 -1950 4487
rect -1916 4453 -1910 4487
rect -2214 4368 -1984 4374
rect -2214 4334 -2115 4368
rect -2081 4334 -2043 4368
rect -2009 4334 -1984 4368
rect -2214 4328 -1984 4334
rect -1956 4328 -1910 4453
rect -1701 4568 -1649 4606
rect -1701 4496 -1649 4516
rect -1701 4406 -1649 4444
rect -1440 4559 -1394 4871
rect -1185 4986 -1133 5024
rect -1185 4914 -1133 4934
rect -1185 4824 -1133 4862
rect -924 4977 -878 5289
rect -669 5404 -617 5442
rect -669 5332 -617 5352
rect -669 5242 -617 5280
rect -408 5395 -362 5707
rect -153 5822 -101 5860
rect -153 5750 -101 5770
rect -153 5660 -101 5698
rect 108 5813 154 6125
rect 363 6240 415 6278
rect 363 6168 415 6188
rect 363 6078 415 6116
rect 624 6231 670 6543
rect 879 6658 931 6696
rect 879 6586 931 6606
rect 879 6496 931 6534
rect 1140 6649 1186 6961
rect 1398 7067 1444 7146
rect 1398 7033 1404 7067
rect 1438 7033 1444 7067
rect 1398 6995 1444 7033
rect 1398 6961 1404 6995
rect 1438 6961 1444 6995
rect 1398 6882 1444 6961
rect 1214 6876 1444 6882
rect 1214 6842 1239 6876
rect 1273 6842 1311 6876
rect 1345 6842 1444 6876
rect 1214 6836 1444 6842
rect 1398 6774 1444 6836
rect 1214 6768 1444 6774
rect 1214 6734 1239 6768
rect 1273 6734 1311 6768
rect 1345 6734 1444 6768
rect 1214 6728 1444 6734
rect 1140 6615 1146 6649
rect 1180 6615 1186 6649
rect 1140 6577 1186 6615
rect 1140 6543 1146 6577
rect 1180 6543 1186 6577
rect 624 6197 630 6231
rect 664 6197 670 6231
rect 624 6159 670 6197
rect 624 6125 630 6159
rect 664 6125 670 6159
rect 108 5779 114 5813
rect 148 5779 154 5813
rect 108 5741 154 5779
rect 108 5707 114 5741
rect 148 5707 154 5741
rect -408 5361 -402 5395
rect -368 5361 -362 5395
rect -408 5323 -362 5361
rect -408 5289 -402 5323
rect -368 5289 -362 5323
rect -924 4943 -918 4977
rect -884 4943 -878 4977
rect -924 4905 -878 4943
rect -924 4871 -918 4905
rect -884 4871 -878 4905
rect -1440 4525 -1434 4559
rect -1400 4525 -1394 4559
rect -1440 4487 -1394 4525
rect -1440 4453 -1434 4487
rect -1400 4453 -1394 4487
rect -2214 4266 -2168 4328
rect -1956 4266 -1468 4269
rect -2214 4260 -1468 4266
rect -2214 4226 -2115 4260
rect -2081 4226 -2043 4260
rect -2009 4226 -1857 4260
rect -1823 4226 -1785 4260
rect -1751 4226 -1599 4260
rect -1565 4226 -1527 4260
rect -1493 4226 -1468 4260
rect -2214 4220 -1468 4226
rect -2214 4141 -2168 4220
rect -2214 4107 -2208 4141
rect -2174 4107 -2168 4141
rect -2214 4069 -2168 4107
rect -2214 4035 -2208 4069
rect -2174 4035 -2168 4069
rect -2214 3956 -2168 4035
rect -1956 4217 -1468 4220
rect -1956 4141 -1910 4217
rect -1956 4107 -1950 4141
rect -1916 4107 -1910 4141
rect -1956 4069 -1910 4107
rect -1956 4035 -1950 4069
rect -1916 4035 -1910 4069
rect -1956 3956 -1910 4035
rect -2214 3950 -1910 3956
rect -2214 3916 -2115 3950
rect -2081 3916 -2043 3950
rect -2009 3916 -1910 3950
rect -2214 3910 -1910 3916
rect -2214 3732 -2168 3910
rect -1956 3732 -1910 3910
rect -1701 4141 -1649 4217
rect -1701 4107 -1692 4141
rect -1658 4107 -1649 4141
rect -1701 4069 -1649 4107
rect -1701 4035 -1692 4069
rect -1658 4035 -1649 4069
rect -1701 3732 -1649 4035
rect -1440 4141 -1394 4453
rect -1185 4568 -1133 4606
rect -1185 4496 -1133 4516
rect -1185 4406 -1133 4444
rect -924 4559 -878 4871
rect -669 4986 -617 5024
rect -669 4914 -617 4934
rect -669 4824 -617 4862
rect -408 4977 -362 5289
rect -153 5404 -101 5442
rect -153 5332 -101 5352
rect -153 5242 -101 5280
rect 108 5395 154 5707
rect 363 5822 415 5860
rect 363 5750 415 5770
rect 363 5660 415 5698
rect 624 5813 670 6125
rect 879 6240 931 6278
rect 879 6168 931 6188
rect 879 6078 931 6116
rect 1140 6231 1186 6543
rect 1398 6649 1444 6728
rect 1398 6615 1404 6649
rect 1438 6615 1444 6649
rect 1398 6577 1444 6615
rect 1398 6543 1404 6577
rect 1438 6543 1444 6577
rect 1398 6464 1444 6543
rect 1214 6458 1444 6464
rect 1214 6424 1239 6458
rect 1273 6424 1311 6458
rect 1345 6424 1444 6458
rect 1214 6418 1444 6424
rect 1398 6356 1444 6418
rect 1214 6350 1444 6356
rect 1214 6316 1239 6350
rect 1273 6316 1311 6350
rect 1345 6316 1444 6350
rect 1214 6310 1444 6316
rect 1140 6197 1146 6231
rect 1180 6197 1186 6231
rect 1140 6159 1186 6197
rect 1140 6125 1146 6159
rect 1180 6125 1186 6159
rect 698 5997 714 6049
rect 766 5997 786 6049
rect 838 5997 872 6049
rect 938 5997 972 6049
rect 1024 5997 1044 6049
rect 1096 5997 1112 6049
rect 698 5889 714 5941
rect 766 5889 786 5941
rect 838 5889 872 5941
rect 938 5889 972 5941
rect 1024 5889 1044 5941
rect 1096 5889 1112 5941
rect 624 5779 630 5813
rect 664 5779 670 5813
rect 624 5741 670 5779
rect 624 5707 630 5741
rect 664 5707 670 5741
rect 182 5579 198 5631
rect 250 5579 270 5631
rect 322 5579 356 5631
rect 422 5579 456 5631
rect 508 5579 528 5631
rect 580 5579 596 5631
rect 182 5471 198 5523
rect 250 5471 270 5523
rect 322 5471 356 5523
rect 422 5471 456 5523
rect 508 5471 528 5523
rect 580 5471 596 5523
rect 108 5361 114 5395
rect 148 5361 154 5395
rect 108 5323 154 5361
rect 108 5289 114 5323
rect 148 5289 154 5323
rect -334 5161 -318 5213
rect -266 5161 -246 5213
rect -194 5161 -160 5213
rect -94 5161 -60 5213
rect -8 5161 12 5213
rect 64 5161 80 5213
rect -334 5053 -318 5105
rect -266 5053 -246 5105
rect -194 5053 -160 5105
rect -94 5053 -60 5105
rect -8 5053 12 5105
rect 64 5053 80 5105
rect -408 4943 -402 4977
rect -368 4943 -362 4977
rect -408 4905 -362 4943
rect -408 4871 -402 4905
rect -368 4871 -362 4905
rect -850 4743 -834 4795
rect -782 4743 -762 4795
rect -710 4743 -676 4795
rect -610 4743 -576 4795
rect -524 4743 -504 4795
rect -452 4743 -436 4795
rect -850 4635 -834 4687
rect -782 4635 -762 4687
rect -710 4635 -676 4687
rect -610 4635 -576 4687
rect -524 4635 -504 4687
rect -452 4635 -436 4687
rect -924 4525 -918 4559
rect -884 4525 -878 4559
rect -924 4487 -878 4525
rect -924 4453 -918 4487
rect -884 4453 -878 4487
rect -1366 4325 -1350 4377
rect -1298 4325 -1278 4377
rect -1226 4325 -1192 4377
rect -1126 4325 -1092 4377
rect -1040 4325 -1020 4377
rect -968 4325 -952 4377
rect -1366 4217 -1350 4269
rect -1298 4217 -1278 4269
rect -1226 4217 -1192 4269
rect -1126 4217 -1092 4269
rect -1040 4217 -1020 4269
rect -968 4217 -952 4269
rect -1440 4107 -1434 4141
rect -1400 4107 -1394 4141
rect -1440 4069 -1394 4107
rect -1440 4035 -1434 4069
rect -1400 4035 -1394 4069
rect -1440 3988 -1394 4035
rect -1185 4150 -1133 4188
rect -1185 4078 -1133 4098
rect -1185 3988 -1133 4026
rect -924 4141 -878 4453
rect -669 4568 -617 4606
rect -669 4496 -617 4516
rect -669 4406 -617 4444
rect -408 4559 -362 4871
rect -153 4986 -101 5024
rect -153 4914 -101 4934
rect -153 4824 -101 4862
rect 108 4977 154 5289
rect 363 5404 415 5442
rect 363 5332 415 5352
rect 363 5242 415 5280
rect 624 5395 670 5707
rect 879 5822 931 5860
rect 879 5750 931 5770
rect 879 5660 931 5698
rect 1140 5813 1186 6125
rect 1398 6231 1444 6310
rect 1398 6197 1404 6231
rect 1438 6197 1444 6231
rect 1398 6159 1444 6197
rect 1398 6125 1404 6159
rect 1438 6125 1444 6159
rect 1398 6046 1444 6125
rect 1214 6040 1444 6046
rect 1214 6006 1239 6040
rect 1273 6006 1311 6040
rect 1345 6006 1444 6040
rect 1214 6000 1444 6006
rect 1398 5938 1444 6000
rect 1214 5932 1444 5938
rect 1214 5898 1239 5932
rect 1273 5898 1311 5932
rect 1345 5898 1444 5932
rect 1214 5892 1444 5898
rect 1140 5779 1146 5813
rect 1180 5779 1186 5813
rect 1140 5741 1186 5779
rect 1140 5707 1146 5741
rect 1180 5707 1186 5741
rect 624 5361 630 5395
rect 664 5361 670 5395
rect 624 5323 670 5361
rect 624 5289 630 5323
rect 664 5289 670 5323
rect 108 4943 114 4977
rect 148 4943 154 4977
rect 108 4905 154 4943
rect 108 4871 114 4905
rect 148 4871 154 4905
rect -408 4525 -402 4559
rect -368 4525 -362 4559
rect -408 4487 -362 4525
rect -408 4453 -402 4487
rect -368 4453 -362 4487
rect -850 4217 -834 4269
rect -782 4217 -762 4269
rect -710 4217 -676 4269
rect -610 4217 -576 4269
rect -524 4217 -504 4269
rect -452 4217 -436 4269
rect -924 4107 -918 4141
rect -884 4107 -878 4141
rect -924 4069 -878 4107
rect -924 4035 -918 4069
rect -884 4035 -878 4069
rect -924 3988 -878 4035
rect -669 4150 -617 4188
rect -669 4078 -617 4098
rect -669 3988 -617 4026
rect -408 4141 -362 4453
rect -153 4568 -101 4606
rect -153 4496 -101 4516
rect -153 4406 -101 4444
rect 108 4559 154 4871
rect 363 4986 415 5024
rect 363 4914 415 4934
rect 363 4824 415 4862
rect 624 4977 670 5289
rect 879 5404 931 5442
rect 879 5332 931 5352
rect 879 5242 931 5280
rect 1140 5395 1186 5707
rect 1398 5813 1444 5892
rect 1398 5779 1404 5813
rect 1438 5779 1444 5813
rect 1398 5741 1444 5779
rect 1398 5707 1404 5741
rect 1438 5707 1444 5741
rect 1398 5628 1444 5707
rect 1214 5622 1444 5628
rect 1214 5588 1239 5622
rect 1273 5588 1311 5622
rect 1345 5588 1444 5622
rect 1214 5582 1444 5588
rect 1398 5520 1444 5582
rect 1214 5514 1444 5520
rect 1214 5480 1239 5514
rect 1273 5480 1311 5514
rect 1345 5480 1444 5514
rect 1214 5474 1444 5480
rect 1140 5361 1146 5395
rect 1180 5361 1186 5395
rect 1140 5323 1186 5361
rect 1140 5289 1146 5323
rect 1180 5289 1186 5323
rect 698 5161 714 5213
rect 766 5161 786 5213
rect 838 5161 872 5213
rect 938 5161 972 5213
rect 1024 5161 1044 5213
rect 1096 5161 1112 5213
rect 698 5053 714 5105
rect 766 5053 786 5105
rect 838 5053 872 5105
rect 938 5053 972 5105
rect 1024 5053 1044 5105
rect 1096 5053 1112 5105
rect 624 4943 630 4977
rect 664 4943 670 4977
rect 624 4905 670 4943
rect 624 4871 630 4905
rect 664 4871 670 4905
rect 182 4743 198 4795
rect 250 4743 270 4795
rect 322 4743 356 4795
rect 422 4743 456 4795
rect 508 4743 528 4795
rect 580 4743 596 4795
rect 182 4635 198 4687
rect 250 4635 270 4687
rect 322 4635 356 4687
rect 422 4635 456 4687
rect 508 4635 528 4687
rect 580 4635 596 4687
rect 108 4525 114 4559
rect 148 4525 154 4559
rect 108 4487 154 4525
rect 108 4453 114 4487
rect 148 4453 154 4487
rect -334 4325 -318 4377
rect -266 4325 -246 4377
rect -194 4325 -160 4377
rect -94 4325 -60 4377
rect -8 4325 12 4377
rect 64 4325 80 4377
rect -334 4217 -318 4269
rect -266 4217 -246 4269
rect -194 4217 -160 4269
rect -94 4217 -60 4269
rect -8 4217 12 4269
rect 64 4217 80 4269
rect -408 4107 -402 4141
rect -368 4107 -362 4141
rect -408 4069 -362 4107
rect -408 4035 -402 4069
rect -368 4035 -362 4069
rect -408 3988 -362 4035
rect -153 4150 -101 4188
rect -153 4078 -101 4098
rect -153 3988 -101 4026
rect 108 4141 154 4453
rect 363 4568 415 4606
rect 363 4496 415 4516
rect 363 4406 415 4444
rect 624 4559 670 4871
rect 879 4986 931 5024
rect 879 4914 931 4934
rect 879 4824 931 4862
rect 1140 4977 1186 5289
rect 1398 5395 1444 5474
rect 1398 5361 1404 5395
rect 1438 5361 1444 5395
rect 1398 5323 1444 5361
rect 1398 5289 1404 5323
rect 1438 5289 1444 5323
rect 1398 5210 1444 5289
rect 1214 5204 1444 5210
rect 1214 5170 1239 5204
rect 1273 5170 1311 5204
rect 1345 5170 1444 5204
rect 1214 5164 1444 5170
rect 1398 5102 1444 5164
rect 1214 5096 1444 5102
rect 1214 5062 1239 5096
rect 1273 5062 1311 5096
rect 1345 5062 1444 5096
rect 1214 5056 1444 5062
rect 1140 4943 1146 4977
rect 1180 4943 1186 4977
rect 1140 4905 1186 4943
rect 1140 4871 1146 4905
rect 1180 4871 1186 4905
rect 1140 4746 1186 4871
rect 1398 4977 1444 5056
rect 1398 4943 1404 4977
rect 1438 4943 1444 4977
rect 1398 4905 1444 4943
rect 1398 4871 1404 4905
rect 1438 4871 1444 4905
rect 1398 4792 1444 4871
rect 1214 4786 1444 4792
rect 1214 4752 1239 4786
rect 1273 4752 1311 4786
rect 1345 4752 1444 4786
rect 1214 4746 1444 4752
rect 698 4684 1186 4687
rect 1398 4684 1444 4746
rect 698 4678 1444 4684
rect 698 4644 723 4678
rect 757 4644 795 4678
rect 829 4644 981 4678
rect 1015 4644 1053 4678
rect 1087 4644 1239 4678
rect 1273 4644 1311 4678
rect 1345 4644 1444 4678
rect 698 4638 1444 4644
rect 698 4635 1186 4638
rect 624 4525 630 4559
rect 664 4525 670 4559
rect 624 4487 670 4525
rect 624 4453 630 4487
rect 664 4453 670 4487
rect 624 4405 670 4453
rect 879 4559 931 4635
rect 879 4525 888 4559
rect 922 4525 931 4559
rect 879 4487 931 4525
rect 879 4453 888 4487
rect 922 4453 931 4487
rect 879 4269 931 4453
rect 1140 4559 1186 4635
rect 1140 4525 1146 4559
rect 1180 4525 1186 4559
rect 1140 4487 1186 4525
rect 1140 4453 1146 4487
rect 1180 4453 1186 4487
rect 1140 4374 1186 4453
rect 1398 4559 1444 4638
rect 1398 4525 1404 4559
rect 1438 4525 1444 4559
rect 1398 4487 1444 4525
rect 1398 4453 1404 4487
rect 1438 4453 1444 4487
rect 1398 4374 1444 4453
rect 1140 4368 1444 4374
rect 1140 4334 1239 4368
rect 1273 4334 1311 4368
rect 1345 4334 1444 4368
rect 1140 4328 1444 4334
rect 1140 4269 1186 4328
rect 182 4260 624 4269
rect 182 4226 207 4260
rect 241 4226 279 4260
rect 313 4226 465 4260
rect 499 4226 537 4260
rect 571 4226 624 4260
rect 182 4217 624 4226
rect 670 4266 1186 4269
rect 1398 4266 1444 4328
rect 670 4260 1444 4266
rect 670 4226 723 4260
rect 757 4226 795 4260
rect 829 4226 981 4260
rect 1015 4226 1053 4260
rect 1087 4226 1239 4260
rect 1273 4226 1311 4260
rect 1345 4226 1444 4260
rect 670 4220 1444 4226
rect 670 4217 1186 4220
rect 108 4107 114 4141
rect 148 4107 154 4141
rect 108 4069 154 4107
rect 108 4035 114 4069
rect 148 4035 154 4069
rect 108 3988 154 4035
rect 363 4141 415 4217
rect 363 4107 372 4141
rect 406 4107 415 4141
rect 363 4069 415 4107
rect 363 4035 372 4069
rect 406 4035 415 4069
rect 363 3732 415 4035
rect 624 4141 670 4188
rect 624 4107 630 4141
rect 664 4107 670 4141
rect 624 4069 670 4107
rect 624 4035 630 4069
rect 664 4035 670 4069
rect 624 3732 670 4035
rect 879 4141 931 4217
rect 879 4107 888 4141
rect 922 4107 931 4141
rect 879 4069 931 4107
rect 879 4035 888 4069
rect 922 4035 931 4069
rect 879 3732 931 4035
rect 1140 4141 1186 4217
rect 1140 4107 1146 4141
rect 1180 4107 1186 4141
rect 1140 4069 1186 4107
rect 1140 4035 1146 4069
rect 1180 4035 1186 4069
rect 1398 4141 1444 4220
rect 1398 4107 1404 4141
rect 1438 4107 1444 4141
rect 1398 4069 1444 4107
rect 1398 4061 1404 4069
rect 1140 3956 1186 4035
rect 1395 4050 1404 4061
rect 1438 4061 1444 4069
rect 3616 7383 3846 7389
rect 3616 7349 3715 7383
rect 3749 7349 3787 7383
rect 3821 7349 3846 7383
rect 3616 7343 3846 7349
rect 3616 7264 3662 7343
rect 3948 7340 3964 7392
rect 4016 7340 4036 7392
rect 4088 7340 4122 7392
rect 4188 7340 4222 7392
rect 4274 7340 4294 7392
rect 4346 7340 4380 7392
rect 4446 7340 4480 7392
rect 4532 7340 4552 7392
rect 4604 7340 4638 7392
rect 4704 7340 4738 7392
rect 4790 7340 4810 7392
rect 4862 7340 4896 7392
rect 4962 7340 4996 7392
rect 5048 7340 5068 7392
rect 5120 7340 5154 7392
rect 5220 7340 5254 7392
rect 5306 7340 5326 7392
rect 5378 7340 5412 7392
rect 5478 7340 5512 7392
rect 5564 7340 5584 7392
rect 5636 7340 5670 7392
rect 5736 7340 5770 7392
rect 5822 7340 5842 7392
rect 5894 7340 5910 7392
rect 6007 7383 6242 7389
rect 6007 7349 6037 7383
rect 6071 7349 6109 7383
rect 6143 7349 6242 7383
rect 6007 7343 6242 7349
rect 3616 7230 3622 7264
rect 3656 7230 3662 7264
rect 3616 7192 3662 7230
rect 3616 7158 3622 7192
rect 3656 7158 3662 7192
rect 3616 7079 3662 7158
rect 3874 7264 3920 7311
rect 3874 7230 3880 7264
rect 3914 7230 3920 7264
rect 3874 7192 3920 7230
rect 3874 7158 3880 7192
rect 3914 7158 3920 7192
rect 3616 7073 3846 7079
rect 3616 7039 3715 7073
rect 3749 7039 3787 7073
rect 3821 7039 3846 7073
rect 3616 7033 3846 7039
rect 3616 6971 3662 7033
rect 3616 6965 3846 6971
rect 3616 6931 3715 6965
rect 3749 6931 3787 6965
rect 3821 6931 3846 6965
rect 3616 6925 3846 6931
rect 3616 6846 3662 6925
rect 3616 6812 3622 6846
rect 3656 6812 3662 6846
rect 3616 6774 3662 6812
rect 3616 6740 3622 6774
rect 3656 6740 3662 6774
rect 3616 6661 3662 6740
rect 3874 6846 3920 7158
rect 4129 7273 4181 7311
rect 4129 7201 4181 7221
rect 4129 7111 4181 7149
rect 4390 7264 4436 7311
rect 4390 7230 4396 7264
rect 4430 7230 4436 7264
rect 4390 7192 4436 7230
rect 4390 7158 4396 7192
rect 4430 7158 4436 7192
rect 3948 6922 3964 6974
rect 4016 6922 4036 6974
rect 4088 6922 4122 6974
rect 4188 6922 4222 6974
rect 4274 6922 4294 6974
rect 4346 6922 4362 6974
rect 3874 6812 3880 6846
rect 3914 6812 3920 6846
rect 3874 6774 3920 6812
rect 3874 6740 3880 6774
rect 3914 6740 3920 6774
rect 3616 6655 3846 6661
rect 3616 6621 3715 6655
rect 3749 6621 3787 6655
rect 3821 6621 3846 6655
rect 3616 6615 3846 6621
rect 3616 6553 3662 6615
rect 3616 6547 3846 6553
rect 3616 6513 3715 6547
rect 3749 6513 3787 6547
rect 3821 6513 3846 6547
rect 3616 6507 3846 6513
rect 3616 6428 3662 6507
rect 3616 6394 3622 6428
rect 3656 6394 3662 6428
rect 3616 6356 3662 6394
rect 3616 6322 3622 6356
rect 3656 6322 3662 6356
rect 3616 6243 3662 6322
rect 3874 6428 3920 6740
rect 4129 6855 4181 6893
rect 4129 6783 4181 6803
rect 4129 6693 4181 6731
rect 4390 6846 4436 7158
rect 4645 7273 4697 7311
rect 4645 7201 4697 7221
rect 4645 7111 4697 7149
rect 4906 7264 4952 7311
rect 4906 7230 4912 7264
rect 4946 7230 4952 7264
rect 4906 7192 4952 7230
rect 4906 7158 4912 7192
rect 4946 7158 4952 7192
rect 4390 6812 4396 6846
rect 4430 6812 4436 6846
rect 4390 6774 4436 6812
rect 4390 6740 4396 6774
rect 4430 6740 4436 6774
rect 3874 6394 3880 6428
rect 3914 6394 3920 6428
rect 3874 6356 3920 6394
rect 3874 6322 3880 6356
rect 3914 6322 3920 6356
rect 3616 6237 3846 6243
rect 3616 6203 3715 6237
rect 3749 6203 3787 6237
rect 3821 6203 3846 6237
rect 3616 6197 3846 6203
rect 3616 6135 3662 6197
rect 3616 6129 3846 6135
rect 3616 6095 3715 6129
rect 3749 6095 3787 6129
rect 3821 6095 3846 6129
rect 3616 6089 3846 6095
rect 3616 6010 3662 6089
rect 3616 5976 3622 6010
rect 3656 5976 3662 6010
rect 3616 5938 3662 5976
rect 3616 5904 3622 5938
rect 3656 5904 3662 5938
rect 3616 5825 3662 5904
rect 3874 6010 3920 6322
rect 4129 6437 4181 6475
rect 4129 6365 4181 6385
rect 4129 6275 4181 6313
rect 4390 6428 4436 6740
rect 4645 6855 4697 6893
rect 4645 6783 4697 6803
rect 4645 6693 4697 6731
rect 4906 6846 4952 7158
rect 5161 7273 5213 7311
rect 5161 7201 5213 7221
rect 5161 7111 5213 7149
rect 5422 7264 5468 7311
rect 5422 7230 5428 7264
rect 5462 7230 5468 7264
rect 5422 7192 5468 7230
rect 5422 7158 5428 7192
rect 5462 7158 5468 7192
rect 4980 6922 4996 6974
rect 5048 6922 5068 6974
rect 5120 6922 5154 6974
rect 5220 6922 5254 6974
rect 5306 6922 5326 6974
rect 5378 6922 5394 6974
rect 4906 6812 4912 6846
rect 4946 6812 4952 6846
rect 4906 6774 4952 6812
rect 4906 6740 4912 6774
rect 4946 6740 4952 6774
rect 4464 6612 4480 6664
rect 4532 6612 4552 6664
rect 4604 6612 4638 6664
rect 4704 6612 4738 6664
rect 4790 6612 4810 6664
rect 4862 6612 4878 6664
rect 4464 6504 4480 6556
rect 4532 6504 4552 6556
rect 4604 6504 4638 6556
rect 4704 6504 4738 6556
rect 4790 6504 4810 6556
rect 4862 6504 4878 6556
rect 4390 6394 4396 6428
rect 4430 6394 4436 6428
rect 4390 6356 4436 6394
rect 4390 6322 4396 6356
rect 4430 6322 4436 6356
rect 3948 6194 3964 6246
rect 4016 6194 4036 6246
rect 4088 6194 4122 6246
rect 4188 6194 4222 6246
rect 4274 6194 4294 6246
rect 4346 6194 4362 6246
rect 3948 6086 3964 6138
rect 4016 6086 4036 6138
rect 4088 6086 4122 6138
rect 4188 6086 4222 6138
rect 4274 6086 4294 6138
rect 4346 6086 4362 6138
rect 3874 5976 3880 6010
rect 3914 5976 3920 6010
rect 3874 5938 3920 5976
rect 3874 5904 3880 5938
rect 3914 5904 3920 5938
rect 3616 5819 3846 5825
rect 3616 5785 3715 5819
rect 3749 5785 3787 5819
rect 3821 5785 3846 5819
rect 3616 5779 3846 5785
rect 3616 5717 3662 5779
rect 3616 5711 3846 5717
rect 3616 5677 3715 5711
rect 3749 5677 3787 5711
rect 3821 5677 3846 5711
rect 3616 5671 3846 5677
rect 3616 5592 3662 5671
rect 3616 5558 3622 5592
rect 3656 5558 3662 5592
rect 3616 5520 3662 5558
rect 3616 5486 3622 5520
rect 3656 5486 3662 5520
rect 3616 5407 3662 5486
rect 3874 5592 3920 5904
rect 4129 6019 4181 6057
rect 4129 5947 4181 5967
rect 4129 5857 4181 5895
rect 4390 6010 4436 6322
rect 4645 6437 4697 6475
rect 4645 6365 4697 6385
rect 4645 6275 4697 6313
rect 4906 6428 4952 6740
rect 5161 6855 5213 6893
rect 5161 6783 5213 6803
rect 5161 6693 5213 6731
rect 5422 6846 5468 7158
rect 5677 7273 5729 7311
rect 5677 7201 5729 7221
rect 5677 7111 5729 7149
rect 5938 7264 5984 7311
rect 5938 7230 5944 7264
rect 5978 7230 5984 7264
rect 5938 7192 5984 7230
rect 5938 7158 5944 7192
rect 5978 7158 5984 7192
rect 5422 6812 5428 6846
rect 5462 6812 5468 6846
rect 5422 6774 5468 6812
rect 5422 6740 5428 6774
rect 5462 6740 5468 6774
rect 4906 6394 4912 6428
rect 4946 6394 4952 6428
rect 4906 6356 4952 6394
rect 4906 6322 4912 6356
rect 4946 6322 4952 6356
rect 4390 5976 4396 6010
rect 4430 5976 4436 6010
rect 4390 5938 4436 5976
rect 4390 5904 4396 5938
rect 4430 5904 4436 5938
rect 3874 5558 3880 5592
rect 3914 5558 3920 5592
rect 3874 5520 3920 5558
rect 3874 5486 3880 5520
rect 3914 5486 3920 5520
rect 3616 5401 3846 5407
rect 3616 5367 3715 5401
rect 3749 5367 3787 5401
rect 3821 5367 3846 5401
rect 3616 5361 3846 5367
rect 3616 5299 3662 5361
rect 3616 5293 3846 5299
rect 3616 5259 3715 5293
rect 3749 5259 3787 5293
rect 3821 5259 3846 5293
rect 3616 5253 3846 5259
rect 3616 5174 3662 5253
rect 3616 5140 3622 5174
rect 3656 5140 3662 5174
rect 3616 5102 3662 5140
rect 3616 5068 3622 5102
rect 3656 5068 3662 5102
rect 3616 4989 3662 5068
rect 3874 5174 3920 5486
rect 4129 5601 4181 5639
rect 4129 5529 4181 5549
rect 4129 5439 4181 5477
rect 4390 5592 4436 5904
rect 4645 6019 4697 6057
rect 4645 5947 4697 5967
rect 4645 5857 4697 5895
rect 4906 6010 4952 6322
rect 5161 6437 5213 6475
rect 5161 6365 5213 6385
rect 5161 6275 5213 6313
rect 5422 6428 5468 6740
rect 5677 6855 5729 6893
rect 5677 6783 5729 6803
rect 5677 6693 5729 6731
rect 5938 6846 5984 7158
rect 6196 7264 6242 7343
rect 6196 7230 6202 7264
rect 6236 7230 6242 7264
rect 6196 7192 6242 7230
rect 6196 7158 6202 7192
rect 6236 7158 6242 7192
rect 6196 7079 6242 7158
rect 6012 7073 6242 7079
rect 6012 7039 6037 7073
rect 6071 7039 6109 7073
rect 6143 7039 6242 7073
rect 6012 7033 6242 7039
rect 6196 6971 6242 7033
rect 6012 6965 6242 6971
rect 6012 6931 6037 6965
rect 6071 6931 6109 6965
rect 6143 6931 6242 6965
rect 6012 6925 6242 6931
rect 5938 6812 5944 6846
rect 5978 6812 5984 6846
rect 5938 6774 5984 6812
rect 5938 6740 5944 6774
rect 5978 6740 5984 6774
rect 5496 6612 5512 6664
rect 5564 6612 5584 6664
rect 5636 6612 5670 6664
rect 5736 6612 5770 6664
rect 5822 6612 5842 6664
rect 5894 6612 5910 6664
rect 5496 6504 5512 6556
rect 5564 6504 5584 6556
rect 5636 6504 5670 6556
rect 5736 6504 5770 6556
rect 5822 6504 5842 6556
rect 5894 6504 5910 6556
rect 5422 6394 5428 6428
rect 5462 6394 5468 6428
rect 5422 6356 5468 6394
rect 5422 6322 5428 6356
rect 5462 6322 5468 6356
rect 4980 6194 4996 6246
rect 5048 6194 5068 6246
rect 5120 6194 5154 6246
rect 5220 6194 5254 6246
rect 5306 6194 5326 6246
rect 5378 6194 5394 6246
rect 4980 6086 4996 6138
rect 5048 6086 5068 6138
rect 5120 6086 5154 6138
rect 5220 6086 5254 6138
rect 5306 6086 5326 6138
rect 5378 6086 5394 6138
rect 4906 5976 4912 6010
rect 4946 5976 4952 6010
rect 4906 5938 4952 5976
rect 4906 5904 4912 5938
rect 4946 5904 4952 5938
rect 4464 5776 4480 5828
rect 4532 5776 4552 5828
rect 4604 5776 4638 5828
rect 4704 5776 4738 5828
rect 4790 5776 4810 5828
rect 4862 5776 4878 5828
rect 4464 5668 4480 5720
rect 4532 5668 4552 5720
rect 4604 5668 4638 5720
rect 4704 5668 4738 5720
rect 4790 5668 4810 5720
rect 4862 5668 4878 5720
rect 4390 5558 4396 5592
rect 4430 5558 4436 5592
rect 4390 5520 4436 5558
rect 4390 5486 4396 5520
rect 4430 5486 4436 5520
rect 3948 5358 3964 5410
rect 4016 5358 4036 5410
rect 4088 5358 4122 5410
rect 4188 5358 4222 5410
rect 4274 5358 4294 5410
rect 4346 5358 4362 5410
rect 3948 5250 3964 5302
rect 4016 5250 4036 5302
rect 4088 5250 4122 5302
rect 4188 5250 4222 5302
rect 4274 5250 4294 5302
rect 4346 5250 4362 5302
rect 3874 5140 3880 5174
rect 3914 5140 3920 5174
rect 3874 5102 3920 5140
rect 3874 5068 3880 5102
rect 3914 5068 3920 5102
rect 3616 4983 3846 4989
rect 3616 4949 3715 4983
rect 3749 4949 3787 4983
rect 3821 4949 3846 4983
rect 3616 4943 3846 4949
rect 3616 4881 3662 4943
rect 3616 4875 3846 4881
rect 3616 4841 3715 4875
rect 3749 4841 3787 4875
rect 3821 4841 3846 4875
rect 3616 4835 3846 4841
rect 3616 4756 3662 4835
rect 3616 4722 3622 4756
rect 3656 4722 3662 4756
rect 3616 4684 3662 4722
rect 3616 4650 3622 4684
rect 3656 4650 3662 4684
rect 3616 4571 3662 4650
rect 3874 4756 3920 5068
rect 4129 5183 4181 5221
rect 4129 5111 4181 5131
rect 4129 5021 4181 5059
rect 4390 5174 4436 5486
rect 4645 5601 4697 5639
rect 4645 5529 4697 5549
rect 4645 5439 4697 5477
rect 4906 5592 4952 5904
rect 5161 6019 5213 6057
rect 5161 5947 5213 5967
rect 5161 5857 5213 5895
rect 5422 6010 5468 6322
rect 5677 6437 5729 6475
rect 5677 6365 5729 6385
rect 5677 6275 5729 6313
rect 5938 6428 5984 6740
rect 6196 6846 6242 6925
rect 6196 6812 6202 6846
rect 6236 6812 6242 6846
rect 6196 6774 6242 6812
rect 6196 6740 6202 6774
rect 6236 6740 6242 6774
rect 6196 6661 6242 6740
rect 6012 6655 6242 6661
rect 6012 6621 6037 6655
rect 6071 6621 6109 6655
rect 6143 6621 6242 6655
rect 6012 6615 6242 6621
rect 6196 6553 6242 6615
rect 6012 6547 6242 6553
rect 6012 6513 6037 6547
rect 6071 6513 6109 6547
rect 6143 6513 6242 6547
rect 6012 6507 6242 6513
rect 5938 6394 5944 6428
rect 5978 6394 5984 6428
rect 5938 6356 5984 6394
rect 5938 6322 5944 6356
rect 5978 6322 5984 6356
rect 5422 5976 5428 6010
rect 5462 5976 5468 6010
rect 5422 5938 5468 5976
rect 5422 5904 5428 5938
rect 5462 5904 5468 5938
rect 4906 5558 4912 5592
rect 4946 5558 4952 5592
rect 4906 5520 4952 5558
rect 4906 5486 4912 5520
rect 4946 5486 4952 5520
rect 4390 5140 4396 5174
rect 4430 5140 4436 5174
rect 4390 5102 4436 5140
rect 4390 5068 4396 5102
rect 4430 5068 4436 5102
rect 3874 4722 3880 4756
rect 3914 4722 3920 4756
rect 3874 4684 3920 4722
rect 3874 4650 3880 4684
rect 3914 4650 3920 4684
rect 3616 4565 3846 4571
rect 3616 4531 3715 4565
rect 3749 4531 3787 4565
rect 3821 4531 3846 4565
rect 3616 4525 3846 4531
rect 3616 4463 3662 4525
rect 3616 4457 3846 4463
rect 3616 4423 3715 4457
rect 3749 4423 3787 4457
rect 3821 4423 3846 4457
rect 3616 4417 3846 4423
rect 3616 4338 3662 4417
rect 3616 4304 3622 4338
rect 3656 4304 3662 4338
rect 3616 4266 3662 4304
rect 3616 4232 3622 4266
rect 3656 4232 3662 4266
rect 3616 4153 3662 4232
rect 3874 4338 3920 4650
rect 4129 4765 4181 4803
rect 4129 4693 4181 4713
rect 4129 4603 4181 4641
rect 4390 4756 4436 5068
rect 4645 5183 4697 5221
rect 4645 5111 4697 5131
rect 4645 5021 4697 5059
rect 4906 5174 4952 5486
rect 5161 5601 5213 5639
rect 5161 5529 5213 5549
rect 5161 5439 5213 5477
rect 5422 5592 5468 5904
rect 5677 6019 5729 6057
rect 5677 5947 5729 5967
rect 5677 5857 5729 5895
rect 5938 6010 5984 6322
rect 6196 6428 6242 6507
rect 6196 6394 6202 6428
rect 6236 6394 6242 6428
rect 6196 6356 6242 6394
rect 6196 6322 6202 6356
rect 6236 6322 6242 6356
rect 6196 6243 6242 6322
rect 6012 6237 6242 6243
rect 6012 6203 6037 6237
rect 6071 6203 6109 6237
rect 6143 6203 6242 6237
rect 6012 6197 6242 6203
rect 6196 6135 6242 6197
rect 6012 6129 6242 6135
rect 6012 6095 6037 6129
rect 6071 6095 6109 6129
rect 6143 6095 6242 6129
rect 6012 6089 6242 6095
rect 5938 5976 5944 6010
rect 5978 5976 5984 6010
rect 5938 5938 5984 5976
rect 5938 5904 5944 5938
rect 5978 5904 5984 5938
rect 5496 5776 5512 5828
rect 5564 5776 5584 5828
rect 5636 5776 5670 5828
rect 5736 5776 5770 5828
rect 5822 5776 5842 5828
rect 5894 5776 5910 5828
rect 5496 5668 5512 5720
rect 5564 5668 5584 5720
rect 5636 5668 5670 5720
rect 5736 5668 5770 5720
rect 5822 5668 5842 5720
rect 5894 5668 5910 5720
rect 5422 5558 5428 5592
rect 5462 5558 5468 5592
rect 5422 5520 5468 5558
rect 5422 5486 5428 5520
rect 5462 5486 5468 5520
rect 4980 5358 4996 5410
rect 5048 5358 5068 5410
rect 5120 5358 5154 5410
rect 5220 5358 5254 5410
rect 5306 5358 5326 5410
rect 5378 5358 5394 5410
rect 4980 5250 4996 5302
rect 5048 5250 5068 5302
rect 5120 5250 5154 5302
rect 5220 5250 5254 5302
rect 5306 5250 5326 5302
rect 5378 5250 5394 5302
rect 4906 5140 4912 5174
rect 4946 5140 4952 5174
rect 4906 5102 4952 5140
rect 4906 5068 4912 5102
rect 4946 5068 4952 5102
rect 4464 4940 4480 4992
rect 4532 4940 4552 4992
rect 4604 4940 4638 4992
rect 4704 4940 4738 4992
rect 4790 4940 4810 4992
rect 4862 4940 4878 4992
rect 4464 4832 4480 4884
rect 4532 4832 4552 4884
rect 4604 4832 4638 4884
rect 4704 4832 4738 4884
rect 4790 4832 4810 4884
rect 4862 4832 4878 4884
rect 4390 4722 4396 4756
rect 4430 4722 4436 4756
rect 4390 4684 4436 4722
rect 4390 4650 4396 4684
rect 4430 4650 4436 4684
rect 3948 4522 3964 4574
rect 4016 4522 4036 4574
rect 4088 4522 4122 4574
rect 4188 4522 4222 4574
rect 4274 4522 4294 4574
rect 4346 4522 4362 4574
rect 3948 4414 3964 4466
rect 4016 4414 4036 4466
rect 4088 4414 4122 4466
rect 4188 4414 4222 4466
rect 4274 4414 4294 4466
rect 4346 4414 4362 4466
rect 3874 4304 3880 4338
rect 3914 4304 3920 4338
rect 3874 4266 3920 4304
rect 3874 4232 3880 4266
rect 3914 4232 3920 4266
rect 3616 4147 3846 4153
rect 3616 4113 3715 4147
rect 3749 4113 3787 4147
rect 3821 4113 3846 4147
rect 3616 4107 3846 4113
rect 1438 4050 1447 4061
rect 1395 3989 1447 3998
rect 1509 4050 1561 4061
rect 1509 3989 1561 3998
rect 1398 3956 1444 3989
rect 1140 3950 1444 3956
rect 1140 3916 1239 3950
rect 1273 3916 1311 3950
rect 1345 3916 1444 3950
rect 1140 3910 1444 3916
rect 1140 3732 1186 3910
rect 1398 3732 1444 3910
rect 3616 3845 3662 4107
rect 3874 3957 3920 4232
rect 4129 4347 4181 4385
rect 4129 4275 4181 4295
rect 4129 4185 4181 4223
rect 4390 4338 4436 4650
rect 4645 4765 4697 4803
rect 4645 4693 4697 4713
rect 4645 4603 4697 4641
rect 4906 4756 4952 5068
rect 5161 5183 5213 5221
rect 5161 5111 5213 5131
rect 5161 5021 5213 5059
rect 5422 5174 5468 5486
rect 5677 5601 5729 5639
rect 5677 5529 5729 5549
rect 5677 5439 5729 5477
rect 5938 5592 5984 5904
rect 6196 6010 6242 6089
rect 6196 5976 6202 6010
rect 6236 5976 6242 6010
rect 6196 5938 6242 5976
rect 6196 5904 6202 5938
rect 6236 5904 6242 5938
rect 6196 5825 6242 5904
rect 6012 5819 6242 5825
rect 6012 5785 6037 5819
rect 6071 5785 6109 5819
rect 6143 5785 6242 5819
rect 6012 5779 6242 5785
rect 6196 5717 6242 5779
rect 6012 5711 6242 5717
rect 6012 5677 6037 5711
rect 6071 5677 6109 5711
rect 6143 5677 6242 5711
rect 6012 5671 6242 5677
rect 5938 5558 5944 5592
rect 5978 5558 5984 5592
rect 5938 5520 5984 5558
rect 5938 5486 5944 5520
rect 5978 5486 5984 5520
rect 5422 5140 5428 5174
rect 5462 5140 5468 5174
rect 5422 5102 5468 5140
rect 5422 5068 5428 5102
rect 5462 5068 5468 5102
rect 4906 4722 4912 4756
rect 4946 4722 4952 4756
rect 4906 4684 4952 4722
rect 4906 4650 4912 4684
rect 4946 4650 4952 4684
rect 4464 4414 4480 4466
rect 4532 4414 4552 4466
rect 4604 4414 4638 4466
rect 4704 4414 4738 4466
rect 4790 4414 4810 4466
rect 4862 4414 4878 4466
rect 4390 4304 4396 4338
rect 4430 4304 4436 4338
rect 4390 4266 4436 4304
rect 4390 4232 4396 4266
rect 4430 4232 4436 4266
rect 4390 3957 4436 4232
rect 4645 4347 4697 4385
rect 4645 4275 4697 4295
rect 4645 4185 4697 4223
rect 4906 4338 4952 4650
rect 5161 4765 5213 4803
rect 5161 4693 5213 4713
rect 5161 4603 5213 4641
rect 5422 4756 5468 5068
rect 5677 5183 5729 5221
rect 5677 5111 5729 5131
rect 5677 5021 5729 5059
rect 5938 5174 5984 5486
rect 6196 5592 6242 5671
rect 6196 5558 6202 5592
rect 6236 5558 6242 5592
rect 6196 5520 6242 5558
rect 6196 5486 6202 5520
rect 6236 5486 6242 5520
rect 6196 5407 6242 5486
rect 6012 5401 6242 5407
rect 6012 5367 6037 5401
rect 6071 5367 6109 5401
rect 6143 5367 6242 5401
rect 6012 5361 6242 5367
rect 6196 5299 6242 5361
rect 6012 5293 6242 5299
rect 6012 5259 6037 5293
rect 6071 5259 6109 5293
rect 6143 5259 6242 5293
rect 6012 5253 6242 5259
rect 5938 5140 5944 5174
rect 5978 5140 5984 5174
rect 5938 5102 5984 5140
rect 5938 5068 5944 5102
rect 5978 5068 5984 5102
rect 5496 4940 5512 4992
rect 5564 4940 5584 4992
rect 5636 4940 5670 4992
rect 5736 4940 5770 4992
rect 5822 4940 5842 4992
rect 5894 4940 5910 4992
rect 5496 4832 5512 4884
rect 5564 4832 5584 4884
rect 5636 4832 5670 4884
rect 5736 4832 5770 4884
rect 5822 4832 5842 4884
rect 5894 4832 5910 4884
rect 5422 4722 5428 4756
rect 5462 4722 5468 4756
rect 5422 4684 5468 4722
rect 5422 4650 5428 4684
rect 5462 4650 5468 4684
rect 4980 4522 4996 4574
rect 5048 4522 5068 4574
rect 5120 4522 5154 4574
rect 5220 4522 5254 4574
rect 5306 4522 5326 4574
rect 5378 4522 5394 4574
rect 4980 4414 4996 4466
rect 5048 4414 5068 4466
rect 5120 4414 5154 4466
rect 5220 4414 5254 4466
rect 5306 4414 5326 4466
rect 5378 4414 5394 4466
rect 4906 4304 4912 4338
rect 4946 4304 4952 4338
rect 4906 4266 4952 4304
rect 4906 4232 4912 4266
rect 4946 4232 4952 4266
rect 4906 3957 4952 4232
rect 5161 4347 5213 4385
rect 5161 4275 5213 4295
rect 5161 4185 5213 4223
rect 5422 4338 5468 4650
rect 5677 4765 5729 4803
rect 5677 4693 5729 4713
rect 5677 4603 5729 4641
rect 5938 4756 5984 5068
rect 6196 5174 6242 5253
rect 6196 5140 6202 5174
rect 6236 5140 6242 5174
rect 6196 5102 6242 5140
rect 6196 5068 6202 5102
rect 6236 5068 6242 5102
rect 6196 4989 6242 5068
rect 6012 4983 6242 4989
rect 6012 4949 6037 4983
rect 6071 4949 6109 4983
rect 6143 4949 6242 4983
rect 6012 4943 6242 4949
rect 6196 4881 6242 4943
rect 6012 4875 6242 4881
rect 6012 4841 6037 4875
rect 6071 4841 6109 4875
rect 6143 4841 6242 4875
rect 6012 4835 6242 4841
rect 5938 4722 5944 4756
rect 5978 4722 5984 4756
rect 5938 4684 5984 4722
rect 5938 4650 5944 4684
rect 5978 4650 5984 4684
rect 5496 4414 5512 4466
rect 5564 4414 5584 4466
rect 5636 4414 5670 4466
rect 5736 4414 5770 4466
rect 5822 4414 5842 4466
rect 5894 4414 5910 4466
rect 5422 4304 5428 4338
rect 5462 4304 5468 4338
rect 5422 4266 5468 4304
rect 5422 4232 5428 4266
rect 5462 4232 5468 4266
rect 5422 3957 5468 4232
rect 5677 4347 5729 4385
rect 5677 4275 5729 4295
rect 5677 4185 5729 4223
rect 5938 4338 5984 4650
rect 6196 4756 6242 4835
rect 6196 4722 6202 4756
rect 6236 4722 6242 4756
rect 6196 4684 6242 4722
rect 6196 4650 6202 4684
rect 6236 4650 6242 4684
rect 6196 4571 6242 4650
rect 6012 4565 6242 4571
rect 6012 4531 6037 4565
rect 6071 4531 6109 4565
rect 6143 4531 6242 4565
rect 6012 4525 6242 4531
rect 6196 4463 6242 4525
rect 6012 4457 6242 4463
rect 6012 4423 6037 4457
rect 6071 4423 6109 4457
rect 6143 4423 6242 4457
rect 6012 4417 6242 4423
rect 5938 4304 5944 4338
rect 5978 4304 5984 4338
rect 5938 4266 5984 4304
rect 5938 4232 5944 4266
rect 5978 4232 5984 4266
rect 5938 3957 5984 4232
rect 6196 4338 6242 4417
rect 6196 4304 6202 4338
rect 6236 4304 6242 4338
rect 6196 4266 6242 4304
rect 6196 4232 6202 4266
rect 6236 4232 6242 4266
rect 6196 4153 6242 4232
rect 6307 4247 6359 4255
rect 6307 4183 6359 4195
rect 6012 4147 6242 4153
rect 6012 4113 6037 4147
rect 6071 4113 6109 4147
rect 6143 4113 6242 4147
rect 6012 4107 6242 4113
rect 3874 3911 5984 3957
rect 6196 4000 6242 4107
rect 6196 3948 6519 4000
rect 6571 3948 6580 4000
rect 6196 3845 6242 3948
rect 3616 3799 6242 3845
rect -2214 3686 1445 3732
rect -2619 3558 -2567 3568
rect -2619 3280 -2567 3506
rect -2619 3216 -2567 3228
rect 7245 3271 7305 7521
rect 9893 7499 9940 7605
rect 10262 7542 10333 7605
rect 10262 7499 10533 7542
rect 9893 7482 10533 7499
rect 9893 7398 10333 7482
rect 8868 7250 9430 7296
rect 8352 6972 8656 6978
rect 8352 6938 8451 6972
rect 8485 6938 8523 6972
rect 8557 6938 8656 6972
rect 8352 6932 8656 6938
rect 8352 6853 8398 6932
rect 8610 6900 8656 6932
rect 8684 6929 8700 6981
rect 8752 6929 8772 6981
rect 8824 6929 8840 6981
rect 8352 6819 8358 6853
rect 8392 6819 8398 6853
rect 8352 6781 8398 6819
rect 8352 6747 8358 6781
rect 8392 6747 8398 6781
rect 8352 6668 8398 6747
rect 8607 6862 8659 6900
rect 8607 6781 8659 6810
rect 8607 6747 8616 6781
rect 8650 6747 8659 6781
rect 8607 6700 8659 6747
rect 8868 6853 8914 7250
rect 8942 6929 8958 6981
rect 9010 6929 9030 6981
rect 9082 6929 9098 6981
rect 9200 6929 9216 6981
rect 9268 6929 9288 6981
rect 9340 6929 9356 6981
rect 8868 6819 8874 6853
rect 8908 6819 8914 6853
rect 8868 6781 8914 6819
rect 8868 6747 8874 6781
rect 8908 6747 8914 6781
rect 8610 6668 8656 6700
rect 8352 6662 8656 6668
rect 8352 6628 8451 6662
rect 8485 6628 8523 6662
rect 8557 6628 8656 6662
rect 8352 6622 8656 6628
rect 8352 6560 8398 6622
rect 8610 6560 8656 6622
rect 8352 6554 8656 6560
rect 8352 6520 8451 6554
rect 8485 6520 8523 6554
rect 8557 6520 8656 6554
rect 8352 6514 8656 6520
rect 8352 6435 8398 6514
rect 8352 6401 8358 6435
rect 8392 6401 8398 6435
rect 8352 6363 8398 6401
rect 8352 6329 8358 6363
rect 8392 6329 8398 6363
rect 8352 6250 8398 6329
rect 8610 6435 8656 6514
rect 8684 6511 8700 6563
rect 8752 6511 8772 6563
rect 8824 6511 8840 6563
rect 8610 6401 8616 6435
rect 8650 6401 8656 6435
rect 8610 6363 8656 6401
rect 8610 6329 8616 6363
rect 8650 6329 8656 6363
rect 8610 6250 8656 6329
rect 8352 6244 8656 6250
rect 8352 6210 8451 6244
rect 8485 6210 8523 6244
rect 8557 6210 8656 6244
rect 8352 6204 8656 6210
rect 8352 6142 8398 6204
rect 8610 6142 8656 6204
rect 8868 6435 8914 6747
rect 9123 6862 9175 6900
rect 9123 6781 9175 6810
rect 9123 6747 9132 6781
rect 9166 6747 9175 6781
rect 9123 6700 9175 6747
rect 9384 6853 9430 7250
rect 9458 6929 9474 6981
rect 9526 6929 9546 6981
rect 9598 6929 9614 6981
rect 9642 6972 9946 6978
rect 9642 6938 9741 6972
rect 9775 6938 9813 6972
rect 9847 6938 9946 6972
rect 9642 6932 9946 6938
rect 9642 6900 9688 6932
rect 9384 6819 9390 6853
rect 9424 6819 9430 6853
rect 9384 6781 9430 6819
rect 9384 6747 9390 6781
rect 9424 6747 9430 6781
rect 8942 6511 8958 6563
rect 9010 6511 9030 6563
rect 9082 6511 9098 6563
rect 8868 6401 8874 6435
rect 8908 6401 8914 6435
rect 8868 6363 8914 6401
rect 8868 6329 8874 6363
rect 8908 6329 8914 6363
rect 8352 6136 8656 6142
rect 8352 6102 8451 6136
rect 8485 6102 8523 6136
rect 8557 6102 8656 6136
rect 8352 6096 8656 6102
rect 8352 6017 8398 6096
rect 8352 5983 8358 6017
rect 8392 5983 8398 6017
rect 8352 5945 8398 5983
rect 8352 5911 8358 5945
rect 8392 5911 8398 5945
rect 8352 5832 8398 5911
rect 8610 6017 8656 6096
rect 8684 6093 8700 6145
rect 8752 6093 8772 6145
rect 8824 6093 8840 6145
rect 8610 5983 8616 6017
rect 8650 5983 8656 6017
rect 8610 5945 8656 5983
rect 8610 5911 8616 5945
rect 8650 5911 8656 5945
rect 8610 5832 8656 5911
rect 8352 5826 8656 5832
rect 8352 5792 8451 5826
rect 8485 5792 8523 5826
rect 8557 5792 8656 5826
rect 8352 5786 8656 5792
rect 8868 6017 8914 6329
rect 9126 6435 9172 6700
rect 9200 6511 9216 6563
rect 9268 6511 9288 6563
rect 9340 6511 9356 6563
rect 9126 6401 9132 6435
rect 9166 6401 9172 6435
rect 9126 6363 9172 6401
rect 9126 6329 9132 6363
rect 9166 6329 9172 6363
rect 8942 6093 8958 6145
rect 9010 6093 9030 6145
rect 9082 6093 9098 6145
rect 8868 5983 8874 6017
rect 8908 5983 8914 6017
rect 8868 5945 8914 5983
rect 8868 5911 8874 5945
rect 8908 5911 8914 5945
rect 8352 5724 8398 5786
rect 8352 5718 8610 5724
rect 8352 5684 8451 5718
rect 8485 5684 8523 5718
rect 8557 5684 8610 5718
rect 8352 5678 8610 5684
rect 8352 5599 8398 5678
rect 8684 5675 8700 5727
rect 8752 5675 8772 5727
rect 8824 5675 8840 5727
rect 8352 5565 8358 5599
rect 8392 5565 8398 5599
rect 8352 5527 8398 5565
rect 8352 5493 8358 5527
rect 8392 5493 8398 5527
rect 8352 5414 8398 5493
rect 8607 5608 8659 5646
rect 8607 5536 8659 5556
rect 8607 5446 8659 5484
rect 8868 5599 8914 5911
rect 9126 6017 9172 6329
rect 9384 6435 9430 6747
rect 9639 6862 9691 6900
rect 9639 6781 9691 6810
rect 9639 6747 9648 6781
rect 9682 6747 9691 6781
rect 9639 6700 9691 6747
rect 9900 6853 9946 6932
rect 9900 6819 9906 6853
rect 9940 6819 9946 6853
rect 9900 6781 9946 6819
rect 9900 6747 9906 6781
rect 9940 6747 9946 6781
rect 9642 6668 9688 6700
rect 9900 6668 9946 6747
rect 9642 6662 9946 6668
rect 9642 6628 9741 6662
rect 9775 6628 9813 6662
rect 9847 6628 9946 6662
rect 9642 6622 9946 6628
rect 9458 6511 9474 6563
rect 9526 6511 9546 6563
rect 9598 6511 9614 6563
rect 9642 6560 9688 6622
rect 9900 6560 9946 6622
rect 9642 6554 9946 6560
rect 9642 6520 9741 6554
rect 9775 6520 9813 6554
rect 9847 6520 9946 6554
rect 9642 6514 9946 6520
rect 9384 6401 9390 6435
rect 9424 6401 9430 6435
rect 9384 6363 9430 6401
rect 9384 6329 9390 6363
rect 9424 6329 9430 6363
rect 9200 6093 9216 6145
rect 9268 6093 9288 6145
rect 9340 6093 9356 6145
rect 9126 5983 9132 6017
rect 9166 5983 9172 6017
rect 9126 5945 9172 5983
rect 9126 5911 9132 5945
rect 9166 5911 9172 5945
rect 9126 5786 9172 5911
rect 9384 6017 9430 6329
rect 9642 6435 9688 6514
rect 9642 6401 9648 6435
rect 9682 6401 9688 6435
rect 9642 6363 9688 6401
rect 9642 6329 9648 6363
rect 9682 6329 9688 6363
rect 9642 6250 9688 6329
rect 9900 6435 9946 6514
rect 9900 6401 9906 6435
rect 9940 6401 9946 6435
rect 9900 6363 9946 6401
rect 9900 6329 9906 6363
rect 9940 6329 9946 6363
rect 9900 6250 9946 6329
rect 9642 6244 9946 6250
rect 9642 6210 9741 6244
rect 9775 6210 9813 6244
rect 9847 6210 9946 6244
rect 9642 6204 9946 6210
rect 9458 6093 9474 6145
rect 9526 6093 9546 6145
rect 9598 6093 9614 6145
rect 9642 6142 9688 6204
rect 9900 6142 9946 6204
rect 9642 6136 9946 6142
rect 9642 6102 9741 6136
rect 9775 6102 9813 6136
rect 9847 6102 9946 6136
rect 9642 6096 9946 6102
rect 9384 5983 9390 6017
rect 9424 5983 9430 6017
rect 9384 5945 9430 5983
rect 9384 5911 9390 5945
rect 9424 5911 9430 5945
rect 8942 5675 8958 5727
rect 9010 5675 9030 5727
rect 9082 5675 9098 5727
rect 9200 5675 9216 5727
rect 9268 5675 9288 5727
rect 9340 5675 9356 5727
rect 8868 5565 8874 5599
rect 8908 5565 8914 5599
rect 8868 5527 8914 5565
rect 8868 5493 8874 5527
rect 8908 5493 8914 5527
rect 8352 5408 8610 5414
rect 8352 5374 8451 5408
rect 8485 5374 8523 5408
rect 8557 5374 8610 5408
rect 8352 5368 8610 5374
rect 8352 5306 8398 5368
rect 8352 5300 8656 5306
rect 8352 5266 8451 5300
rect 8485 5266 8523 5300
rect 8557 5266 8656 5300
rect 8352 5260 8656 5266
rect 8352 5181 8398 5260
rect 8352 5147 8358 5181
rect 8392 5147 8398 5181
rect 8352 5109 8398 5147
rect 8352 5075 8358 5109
rect 8392 5075 8398 5109
rect 8352 4996 8398 5075
rect 8610 5181 8656 5260
rect 8684 5257 8700 5309
rect 8752 5257 8772 5309
rect 8824 5257 8840 5309
rect 8610 5147 8616 5181
rect 8650 5147 8656 5181
rect 8610 5109 8656 5147
rect 8610 5075 8616 5109
rect 8650 5075 8656 5109
rect 8610 4996 8656 5075
rect 8352 4990 8656 4996
rect 8352 4956 8451 4990
rect 8485 4956 8523 4990
rect 8557 4956 8656 4990
rect 8352 4950 8656 4956
rect 8352 4888 8398 4950
rect 8610 4888 8656 4950
rect 8868 5181 8914 5493
rect 9123 5608 9175 5646
rect 9123 5536 9175 5556
rect 9123 5446 9175 5484
rect 9384 5599 9430 5911
rect 9642 6017 9688 6096
rect 9642 5983 9648 6017
rect 9682 5983 9688 6017
rect 9642 5945 9688 5983
rect 9642 5911 9648 5945
rect 9682 5911 9688 5945
rect 9642 5832 9688 5911
rect 9900 6017 9946 6096
rect 9900 5983 9906 6017
rect 9940 5983 9946 6017
rect 9900 5945 9946 5983
rect 9900 5911 9906 5945
rect 9940 5911 9946 5945
rect 9900 5832 9946 5911
rect 9642 5826 9946 5832
rect 9642 5792 9741 5826
rect 9775 5792 9813 5826
rect 9847 5792 9946 5826
rect 9642 5786 9946 5792
rect 9458 5675 9474 5727
rect 9526 5675 9546 5727
rect 9598 5675 9614 5727
rect 9900 5724 9946 5786
rect 9688 5718 9946 5724
rect 9688 5684 9741 5718
rect 9775 5684 9813 5718
rect 9847 5684 9946 5718
rect 9688 5678 9946 5684
rect 9384 5565 9390 5599
rect 9424 5565 9430 5599
rect 9384 5527 9430 5565
rect 9384 5493 9390 5527
rect 9424 5493 9430 5527
rect 8942 5257 8958 5309
rect 9010 5257 9030 5309
rect 9082 5257 9098 5309
rect 8868 5147 8874 5181
rect 8908 5147 8914 5181
rect 8868 5109 8914 5147
rect 8868 5075 8874 5109
rect 8908 5075 8914 5109
rect 8352 4882 8656 4888
rect 8352 4848 8451 4882
rect 8485 4848 8523 4882
rect 8557 4848 8656 4882
rect 8352 4842 8656 4848
rect 8352 4763 8398 4842
rect 8352 4729 8358 4763
rect 8392 4729 8398 4763
rect 8352 4691 8398 4729
rect 8352 4657 8358 4691
rect 8392 4657 8398 4691
rect 8352 4578 8398 4657
rect 8610 4763 8656 4842
rect 8684 4839 8700 4891
rect 8752 4839 8772 4891
rect 8824 4839 8840 4891
rect 8610 4729 8616 4763
rect 8650 4729 8656 4763
rect 8610 4691 8656 4729
rect 8610 4657 8616 4691
rect 8650 4657 8656 4691
rect 8610 4578 8656 4657
rect 8352 4572 8656 4578
rect 8352 4538 8451 4572
rect 8485 4538 8523 4572
rect 8557 4538 8656 4572
rect 8352 4532 8656 4538
rect 8352 4470 8398 4532
rect 8610 4470 8656 4532
rect 8868 4763 8914 5075
rect 9126 5181 9172 5306
rect 9200 5257 9216 5309
rect 9268 5257 9288 5309
rect 9340 5257 9356 5309
rect 9126 5147 9132 5181
rect 9166 5147 9172 5181
rect 9126 5109 9172 5147
rect 9126 5075 9132 5109
rect 9166 5075 9172 5109
rect 8942 4839 8958 4891
rect 9010 4839 9030 4891
rect 9082 4839 9098 4891
rect 8868 4729 8874 4763
rect 8908 4729 8914 4763
rect 8868 4691 8914 4729
rect 8868 4657 8874 4691
rect 8908 4657 8914 4691
rect 8352 4464 8656 4470
rect 8352 4430 8451 4464
rect 8485 4430 8523 4464
rect 8557 4430 8656 4464
rect 8352 4424 8656 4430
rect 8352 4345 8398 4424
rect 8352 4311 8358 4345
rect 8392 4311 8398 4345
rect 8352 4273 8398 4311
rect 8352 4239 8358 4273
rect 8392 4239 8398 4273
rect 8352 4160 8398 4239
rect 8610 4345 8656 4424
rect 8684 4421 8700 4473
rect 8752 4421 8772 4473
rect 8824 4421 8840 4473
rect 8610 4311 8616 4345
rect 8650 4311 8656 4345
rect 8610 4273 8656 4311
rect 8610 4239 8616 4273
rect 8650 4239 8656 4273
rect 8610 4160 8656 4239
rect 8868 4345 8914 4657
rect 9126 4763 9172 5075
rect 9384 5181 9430 5493
rect 9639 5608 9691 5646
rect 9639 5536 9691 5556
rect 9639 5446 9691 5484
rect 9900 5599 9946 5678
rect 9900 5565 9906 5599
rect 9940 5565 9946 5599
rect 9900 5527 9946 5565
rect 9900 5493 9906 5527
rect 9940 5493 9946 5527
rect 9900 5414 9946 5493
rect 9688 5408 9946 5414
rect 9688 5374 9741 5408
rect 9775 5374 9813 5408
rect 9847 5374 9946 5408
rect 9688 5368 9946 5374
rect 9458 5257 9474 5309
rect 9526 5257 9546 5309
rect 9598 5257 9614 5309
rect 9900 5306 9946 5368
rect 9642 5300 9946 5306
rect 9642 5266 9741 5300
rect 9775 5266 9813 5300
rect 9847 5266 9946 5300
rect 9642 5260 9946 5266
rect 9384 5147 9390 5181
rect 9424 5147 9430 5181
rect 9384 5109 9430 5147
rect 9384 5075 9390 5109
rect 9424 5075 9430 5109
rect 9200 4839 9216 4891
rect 9268 4839 9288 4891
rect 9340 4839 9356 4891
rect 9126 4729 9132 4763
rect 9166 4729 9172 4763
rect 9126 4691 9172 4729
rect 9126 4657 9132 4691
rect 9166 4657 9172 4691
rect 8942 4421 8958 4473
rect 9010 4421 9030 4473
rect 9082 4421 9098 4473
rect 8868 4311 8874 4345
rect 8908 4311 8914 4345
rect 8868 4273 8914 4311
rect 8868 4239 8874 4273
rect 8908 4239 8914 4273
rect 8868 4192 8914 4239
rect 9126 4345 9172 4657
rect 9384 4763 9430 5075
rect 9642 5181 9688 5260
rect 9642 5147 9648 5181
rect 9682 5147 9688 5181
rect 9642 5109 9688 5147
rect 9642 5075 9648 5109
rect 9682 5075 9688 5109
rect 9642 4996 9688 5075
rect 9900 5181 9946 5260
rect 9900 5147 9906 5181
rect 9940 5147 9946 5181
rect 9900 5109 9946 5147
rect 9900 5075 9906 5109
rect 9940 5075 9946 5109
rect 9900 4996 9946 5075
rect 9642 4990 9946 4996
rect 9642 4956 9741 4990
rect 9775 4956 9813 4990
rect 9847 4956 9946 4990
rect 9642 4950 9946 4956
rect 9458 4839 9474 4891
rect 9526 4839 9546 4891
rect 9598 4839 9614 4891
rect 9642 4888 9688 4950
rect 9900 4888 9946 4950
rect 9642 4882 9946 4888
rect 9642 4848 9741 4882
rect 9775 4848 9813 4882
rect 9847 4848 9946 4882
rect 9642 4842 9946 4848
rect 9384 4729 9390 4763
rect 9424 4729 9430 4763
rect 9384 4691 9430 4729
rect 9384 4657 9390 4691
rect 9424 4657 9430 4691
rect 9200 4421 9216 4473
rect 9268 4421 9288 4473
rect 9340 4421 9356 4473
rect 9126 4311 9132 4345
rect 9166 4311 9172 4345
rect 9126 4273 9172 4311
rect 9126 4239 9132 4273
rect 9166 4239 9172 4273
rect 8352 4154 8656 4160
rect 8352 4120 8451 4154
rect 8485 4120 8523 4154
rect 8557 4120 8656 4154
rect 8352 4114 8656 4120
rect 8352 3808 8398 4114
rect 8335 3796 8415 3808
rect 8335 3744 8349 3796
rect 8401 3744 8415 3796
rect 8335 3732 8415 3744
rect 8610 3732 8656 4114
rect 9126 3732 9172 4239
rect 9384 4345 9430 4657
rect 9642 4763 9688 4842
rect 9642 4729 9648 4763
rect 9682 4729 9688 4763
rect 9642 4691 9688 4729
rect 9642 4657 9648 4691
rect 9682 4657 9688 4691
rect 9642 4578 9688 4657
rect 9900 4763 9946 4842
rect 9900 4729 9906 4763
rect 9940 4729 9946 4763
rect 9900 4691 9946 4729
rect 9900 4657 9906 4691
rect 9940 4657 9946 4691
rect 9900 4578 9946 4657
rect 9642 4572 9946 4578
rect 9642 4538 9741 4572
rect 9775 4538 9813 4572
rect 9847 4538 9946 4572
rect 9642 4532 9946 4538
rect 9458 4421 9474 4473
rect 9526 4421 9546 4473
rect 9598 4421 9614 4473
rect 9642 4470 9688 4532
rect 9900 4470 9946 4532
rect 9642 4464 9946 4470
rect 9642 4430 9741 4464
rect 9775 4430 9813 4464
rect 9847 4430 9946 4464
rect 9642 4424 9946 4430
rect 9384 4311 9390 4345
rect 9424 4311 9430 4345
rect 9384 4273 9430 4311
rect 9384 4239 9390 4273
rect 9424 4239 9430 4273
rect 9384 4192 9430 4239
rect 9642 4345 9688 4424
rect 9642 4311 9648 4345
rect 9682 4311 9688 4345
rect 9642 4273 9688 4311
rect 9642 4239 9648 4273
rect 9682 4239 9688 4273
rect 9642 4160 9688 4239
rect 9900 4345 9946 4424
rect 9900 4311 9906 4345
rect 9940 4311 9946 4345
rect 9900 4273 9946 4311
rect 9900 4239 9906 4273
rect 9940 4239 9946 4273
rect 9900 4160 9946 4239
rect 9642 4154 9946 4160
rect 9642 4120 9741 4154
rect 9775 4120 9813 4154
rect 9847 4120 9946 4154
rect 9642 4114 9946 4120
rect 9642 3732 9688 4114
rect 9900 4052 9946 4114
rect 9900 4018 9906 4052
rect 9940 4018 9946 4052
rect 9900 3732 9946 4018
rect 10487 3732 10533 7482
rect 11103 4292 11163 8004
rect 11062 4247 11214 4292
rect 11062 4195 11107 4247
rect 11159 4195 11214 4247
rect 11062 4148 11214 4195
rect 8352 3686 10533 3732
rect 7245 3219 7249 3271
rect 7301 3219 7305 3271
rect 7245 3192 7305 3219
<< via1 >>
rect -897 10233 -845 10242
rect -897 10199 -888 10233
rect -888 10199 -854 10233
rect -854 10199 -845 10233
rect -897 10190 -845 10199
rect -825 10233 -773 10242
rect -825 10199 -816 10233
rect -816 10199 -782 10233
rect -782 10199 -773 10233
rect -825 10190 -773 10199
rect -639 10233 -587 10242
rect -639 10199 -630 10233
rect -630 10199 -596 10233
rect -596 10199 -587 10233
rect -639 10190 -587 10199
rect -567 10233 -515 10242
rect -567 10199 -558 10233
rect -558 10199 -524 10233
rect -524 10199 -515 10233
rect -567 10190 -515 10199
rect -897 10125 -845 10134
rect -897 10091 -888 10125
rect -888 10091 -854 10125
rect -854 10091 -845 10125
rect -897 10082 -845 10091
rect -825 10125 -773 10134
rect -825 10091 -816 10125
rect -816 10091 -782 10125
rect -782 10091 -773 10125
rect -825 10082 -773 10091
rect -639 10125 -587 10134
rect -639 10091 -630 10125
rect -630 10091 -596 10125
rect -596 10091 -587 10125
rect -639 10082 -587 10091
rect -567 10125 -515 10134
rect -567 10091 -558 10125
rect -558 10091 -524 10125
rect -524 10091 -515 10125
rect -567 10082 -515 10091
rect -732 9997 -680 10006
rect -732 9963 -723 9997
rect -723 9963 -689 9997
rect -689 9963 -680 9997
rect -732 9954 -680 9963
rect -732 9925 -680 9934
rect -732 9891 -723 9925
rect -723 9891 -689 9925
rect -689 9891 -680 9925
rect -732 9882 -680 9891
rect -216 10433 -164 10442
rect -216 10399 -207 10433
rect -207 10399 -173 10433
rect -173 10399 -164 10433
rect -216 10390 -164 10399
rect -216 10361 -164 10370
rect -216 10327 -207 10361
rect -207 10327 -173 10361
rect -173 10327 -164 10361
rect -216 10318 -164 10327
rect -381 10233 -329 10242
rect -381 10199 -372 10233
rect -372 10199 -338 10233
rect -338 10199 -329 10233
rect -381 10190 -329 10199
rect -309 10233 -257 10242
rect -309 10199 -300 10233
rect -300 10199 -266 10233
rect -266 10199 -257 10233
rect -309 10190 -257 10199
rect -123 10233 -71 10242
rect -123 10199 -114 10233
rect -114 10199 -80 10233
rect -80 10199 -71 10233
rect -123 10190 -71 10199
rect -51 10233 1 10242
rect -51 10199 -42 10233
rect -42 10199 -8 10233
rect -8 10199 1 10233
rect -51 10190 1 10199
rect -381 10125 -329 10134
rect -381 10091 -372 10125
rect -372 10091 -338 10125
rect -338 10091 -329 10125
rect -381 10082 -329 10091
rect -309 10125 -257 10134
rect -309 10091 -300 10125
rect -300 10091 -266 10125
rect -266 10091 -257 10125
rect -309 10082 -257 10091
rect -123 10125 -71 10134
rect -123 10091 -114 10125
rect -114 10091 -80 10125
rect -80 10091 -71 10125
rect -123 10082 -71 10091
rect -51 10125 1 10134
rect -51 10091 -42 10125
rect -42 10091 -8 10125
rect -8 10091 1 10125
rect -51 10082 1 10091
rect -897 9361 -845 9370
rect -897 9327 -888 9361
rect -888 9327 -854 9361
rect -854 9327 -845 9361
rect -897 9318 -845 9327
rect -825 9361 -773 9370
rect -825 9327 -816 9361
rect -816 9327 -782 9361
rect -782 9327 -773 9361
rect -825 9318 -773 9327
rect -639 9361 -587 9370
rect -639 9327 -630 9361
rect -630 9327 -596 9361
rect -596 9327 -587 9361
rect -639 9318 -587 9327
rect -567 9361 -515 9370
rect -567 9327 -558 9361
rect -558 9327 -524 9361
rect -524 9327 -515 9361
rect -567 9318 -515 9327
rect -897 9253 -845 9262
rect -897 9219 -888 9253
rect -888 9219 -854 9253
rect -854 9219 -845 9253
rect -897 9210 -845 9219
rect -825 9253 -773 9262
rect -825 9219 -816 9253
rect -816 9219 -782 9253
rect -782 9219 -773 9253
rect -825 9210 -773 9219
rect -639 9253 -587 9262
rect -639 9219 -630 9253
rect -630 9219 -596 9253
rect -596 9219 -587 9253
rect -639 9210 -587 9219
rect -567 9253 -515 9262
rect -567 9219 -558 9253
rect -558 9219 -524 9253
rect -524 9219 -515 9253
rect -567 9210 -515 9219
rect -732 9125 -680 9134
rect -732 9091 -723 9125
rect -723 9091 -689 9125
rect -689 9091 -680 9125
rect -732 9082 -680 9091
rect -732 9053 -680 9062
rect -732 9019 -723 9053
rect -723 9019 -689 9053
rect -689 9019 -680 9053
rect -732 9010 -680 9019
rect -216 9561 -164 9570
rect -216 9527 -207 9561
rect -207 9527 -173 9561
rect -173 9527 -164 9561
rect -216 9518 -164 9527
rect -216 9489 -164 9498
rect -216 9455 -207 9489
rect -207 9455 -173 9489
rect -173 9455 -164 9489
rect -216 9446 -164 9455
rect -381 9361 -329 9370
rect -381 9327 -372 9361
rect -372 9327 -338 9361
rect -338 9327 -329 9361
rect -381 9318 -329 9327
rect -309 9361 -257 9370
rect -309 9327 -300 9361
rect -300 9327 -266 9361
rect -266 9327 -257 9361
rect -309 9318 -257 9327
rect -123 9361 -71 9370
rect -123 9327 -114 9361
rect -114 9327 -80 9361
rect -80 9327 -71 9361
rect -123 9318 -71 9327
rect -51 9361 1 9370
rect -51 9327 -42 9361
rect -42 9327 -8 9361
rect -8 9327 1 9361
rect -51 9318 1 9327
rect -381 9253 -329 9262
rect -381 9219 -372 9253
rect -372 9219 -338 9253
rect -338 9219 -329 9253
rect -381 9210 -329 9219
rect -309 9253 -257 9262
rect -309 9219 -300 9253
rect -300 9219 -266 9253
rect -266 9219 -257 9253
rect -309 9210 -257 9219
rect -123 9253 -71 9262
rect -123 9219 -114 9253
rect -114 9219 -80 9253
rect -80 9219 -71 9253
rect -123 9210 -71 9219
rect -51 9253 1 9262
rect -51 9219 -42 9253
rect -42 9219 -8 9253
rect -8 9219 1 9253
rect -51 9210 1 9219
rect 3683 10771 3735 10780
rect 3683 10737 3692 10771
rect 3692 10737 3726 10771
rect 3726 10737 3735 10771
rect 3683 10728 3735 10737
rect 3755 10771 3807 10780
rect 3755 10737 3764 10771
rect 3764 10737 3798 10771
rect 3798 10737 3807 10771
rect 3755 10728 3807 10737
rect 4457 10771 4509 10780
rect 4457 10737 4466 10771
rect 4466 10737 4500 10771
rect 4500 10737 4509 10771
rect 4457 10728 4509 10737
rect 4529 10771 4581 10780
rect 4529 10737 4538 10771
rect 4538 10737 4572 10771
rect 4572 10737 4581 10771
rect 4529 10728 4581 10737
rect 3590 10652 3642 10661
rect 3590 10618 3599 10652
rect 3599 10618 3633 10652
rect 3633 10618 3642 10652
rect 3590 10609 3642 10618
rect 3590 10580 3642 10589
rect 3590 10546 3599 10580
rect 3599 10546 3633 10580
rect 3633 10546 3642 10580
rect 3590 10537 3642 10546
rect 3590 10234 3642 10243
rect 3590 10200 3599 10234
rect 3599 10200 3633 10234
rect 3633 10200 3642 10234
rect 3590 10191 3642 10200
rect 3590 10162 3642 10171
rect 3590 10128 3599 10162
rect 3599 10128 3633 10162
rect 3633 10128 3642 10162
rect 3590 10119 3642 10128
rect 4106 10652 4158 10661
rect 4106 10618 4115 10652
rect 4115 10618 4149 10652
rect 4149 10618 4158 10652
rect 4106 10609 4158 10618
rect 4106 10580 4158 10589
rect 4106 10546 4115 10580
rect 4115 10546 4149 10580
rect 4149 10546 4158 10580
rect 4106 10537 4158 10546
rect 3941 10461 3993 10467
rect 3941 10427 3950 10461
rect 3950 10427 3984 10461
rect 3984 10427 3993 10461
rect 3941 10415 3993 10427
rect 4013 10461 4065 10467
rect 4013 10427 4022 10461
rect 4022 10427 4056 10461
rect 4056 10427 4065 10461
rect 4013 10415 4065 10427
rect 4199 10461 4251 10467
rect 4199 10427 4208 10461
rect 4208 10427 4242 10461
rect 4242 10427 4251 10461
rect 4199 10415 4251 10427
rect 4271 10461 4323 10467
rect 4271 10427 4280 10461
rect 4280 10427 4314 10461
rect 4314 10427 4323 10461
rect 4271 10415 4323 10427
rect 3941 10353 3993 10362
rect 3941 10319 3950 10353
rect 3950 10319 3984 10353
rect 3984 10319 3993 10353
rect 3941 10310 3993 10319
rect 4013 10353 4065 10362
rect 4013 10319 4022 10353
rect 4022 10319 4056 10353
rect 4056 10319 4065 10353
rect 4013 10310 4065 10319
rect 4199 10353 4251 10362
rect 4199 10319 4208 10353
rect 4208 10319 4242 10353
rect 4242 10319 4251 10353
rect 4199 10310 4251 10319
rect 4271 10353 4323 10362
rect 4271 10319 4280 10353
rect 4280 10319 4314 10353
rect 4314 10319 4323 10353
rect 4271 10310 4323 10319
rect 3425 10043 3477 10049
rect 3425 10009 3434 10043
rect 3434 10009 3468 10043
rect 3468 10009 3477 10043
rect 3425 9997 3477 10009
rect 3497 10043 3549 10049
rect 3497 10009 3506 10043
rect 3506 10009 3540 10043
rect 3540 10009 3549 10043
rect 3497 9997 3549 10009
rect 3683 10043 3735 10049
rect 3683 10009 3692 10043
rect 3692 10009 3726 10043
rect 3726 10009 3735 10043
rect 3683 9997 3735 10009
rect 3755 10043 3807 10049
rect 3755 10009 3764 10043
rect 3764 10009 3798 10043
rect 3798 10009 3807 10043
rect 3755 9997 3807 10009
rect 3425 9935 3477 9944
rect 3425 9901 3434 9935
rect 3434 9901 3468 9935
rect 3468 9901 3477 9935
rect 3425 9892 3477 9901
rect 3497 9935 3549 9944
rect 3497 9901 3506 9935
rect 3506 9901 3540 9935
rect 3540 9901 3549 9935
rect 3497 9892 3549 9901
rect 3683 9935 3735 9944
rect 3683 9901 3692 9935
rect 3692 9901 3726 9935
rect 3726 9901 3735 9935
rect 3683 9892 3735 9901
rect 3755 9935 3807 9944
rect 3755 9901 3764 9935
rect 3764 9901 3798 9935
rect 3798 9901 3807 9935
rect 3755 9892 3807 9901
rect 3590 9816 3642 9825
rect 3590 9782 3599 9816
rect 3599 9782 3633 9816
rect 3633 9782 3642 9816
rect 3590 9773 3642 9782
rect 3590 9744 3642 9753
rect 3590 9710 3599 9744
rect 3599 9710 3633 9744
rect 3633 9710 3642 9744
rect 3590 9701 3642 9710
rect 4106 10234 4158 10243
rect 4106 10200 4115 10234
rect 4115 10200 4149 10234
rect 4149 10200 4158 10234
rect 4106 10191 4158 10200
rect 4106 10162 4158 10171
rect 4106 10128 4115 10162
rect 4115 10128 4149 10162
rect 4149 10128 4158 10162
rect 4106 10119 4158 10128
rect 4622 10652 4674 10661
rect 4622 10618 4631 10652
rect 4631 10618 4665 10652
rect 4665 10618 4674 10652
rect 4622 10609 4674 10618
rect 4622 10580 4674 10589
rect 4622 10546 4631 10580
rect 4631 10546 4665 10580
rect 4665 10546 4674 10580
rect 4622 10537 4674 10546
rect 3590 9398 3642 9407
rect 3590 9364 3599 9398
rect 3599 9364 3633 9398
rect 3633 9364 3642 9398
rect 3590 9355 3642 9364
rect 3590 9326 3642 9335
rect 3590 9292 3599 9326
rect 3599 9292 3633 9326
rect 3633 9292 3642 9326
rect 3590 9283 3642 9292
rect 4106 9816 4158 9825
rect 4106 9782 4115 9816
rect 4115 9782 4149 9816
rect 4149 9782 4158 9816
rect 4106 9773 4158 9782
rect 4106 9744 4158 9753
rect 4106 9710 4115 9744
rect 4115 9710 4149 9744
rect 4149 9710 4158 9744
rect 4106 9701 4158 9710
rect 4622 10234 4674 10243
rect 4622 10200 4631 10234
rect 4631 10200 4665 10234
rect 4665 10200 4674 10234
rect 4622 10191 4674 10200
rect 4622 10162 4674 10171
rect 4622 10128 4631 10162
rect 4631 10128 4665 10162
rect 4665 10128 4674 10162
rect 4622 10119 4674 10128
rect 4457 10043 4509 10049
rect 4457 10009 4466 10043
rect 4466 10009 4500 10043
rect 4500 10009 4509 10043
rect 4457 9997 4509 10009
rect 4529 10043 4581 10049
rect 4529 10009 4538 10043
rect 4538 10009 4572 10043
rect 4572 10009 4581 10043
rect 4529 9997 4581 10009
rect 4715 10043 4767 10049
rect 4715 10009 4724 10043
rect 4724 10009 4758 10043
rect 4758 10009 4767 10043
rect 4715 9997 4767 10009
rect 4787 10043 4839 10049
rect 4787 10009 4796 10043
rect 4796 10009 4830 10043
rect 4830 10009 4839 10043
rect 4787 9997 4839 10009
rect 4457 9935 4509 9944
rect 4457 9901 4466 9935
rect 4466 9901 4500 9935
rect 4500 9901 4509 9935
rect 4457 9892 4509 9901
rect 4529 9935 4581 9944
rect 4529 9901 4538 9935
rect 4538 9901 4572 9935
rect 4572 9901 4581 9935
rect 4529 9892 4581 9901
rect 4715 9935 4767 9944
rect 4715 9901 4724 9935
rect 4724 9901 4758 9935
rect 4758 9901 4767 9935
rect 4715 9892 4767 9901
rect 4787 9935 4839 9944
rect 4787 9901 4796 9935
rect 4796 9901 4830 9935
rect 4830 9901 4839 9935
rect 4787 9892 4839 9901
rect 3941 9625 3993 9631
rect 3941 9591 3950 9625
rect 3950 9591 3984 9625
rect 3984 9591 3993 9625
rect 3941 9579 3993 9591
rect 4013 9625 4065 9631
rect 4013 9591 4022 9625
rect 4022 9591 4056 9625
rect 4056 9591 4065 9625
rect 4013 9579 4065 9591
rect 4199 9625 4251 9631
rect 4199 9591 4208 9625
rect 4208 9591 4242 9625
rect 4242 9591 4251 9625
rect 4199 9579 4251 9591
rect 4271 9625 4323 9631
rect 4271 9591 4280 9625
rect 4280 9591 4314 9625
rect 4314 9591 4323 9625
rect 4271 9579 4323 9591
rect 3941 9517 3993 9526
rect 3941 9483 3950 9517
rect 3950 9483 3984 9517
rect 3984 9483 3993 9517
rect 3941 9474 3993 9483
rect 4013 9517 4065 9526
rect 4013 9483 4022 9517
rect 4022 9483 4056 9517
rect 4056 9483 4065 9517
rect 4013 9474 4065 9483
rect 4199 9517 4251 9526
rect 4199 9483 4208 9517
rect 4208 9483 4242 9517
rect 4242 9483 4251 9517
rect 4199 9474 4251 9483
rect 4271 9517 4323 9526
rect 4271 9483 4280 9517
rect 4280 9483 4314 9517
rect 4314 9483 4323 9517
rect 4271 9474 4323 9483
rect 3425 9207 3477 9213
rect 3425 9173 3434 9207
rect 3434 9173 3468 9207
rect 3468 9173 3477 9207
rect 3425 9161 3477 9173
rect 3497 9207 3549 9213
rect 3497 9173 3506 9207
rect 3506 9173 3540 9207
rect 3540 9173 3549 9207
rect 3497 9161 3549 9173
rect 3683 9207 3735 9213
rect 3683 9173 3692 9207
rect 3692 9173 3726 9207
rect 3726 9173 3735 9207
rect 3683 9161 3735 9173
rect 3755 9207 3807 9213
rect 3755 9173 3764 9207
rect 3764 9173 3798 9207
rect 3798 9173 3807 9207
rect 3755 9161 3807 9173
rect 3425 9095 3477 9104
rect 3425 9061 3434 9095
rect 3434 9061 3468 9095
rect 3468 9061 3477 9095
rect 3425 9052 3477 9061
rect 3497 9095 3549 9104
rect 3497 9061 3506 9095
rect 3506 9061 3540 9095
rect 3540 9061 3549 9095
rect 3497 9052 3549 9061
rect 3683 9095 3735 9104
rect 3683 9061 3692 9095
rect 3692 9061 3726 9095
rect 3726 9061 3735 9095
rect 3683 9052 3735 9061
rect 3755 9095 3807 9104
rect 3755 9061 3764 9095
rect 3764 9061 3798 9095
rect 3798 9061 3807 9095
rect 3755 9052 3807 9061
rect 3590 8976 3642 8985
rect 3590 8942 3599 8976
rect 3599 8942 3633 8976
rect 3633 8942 3642 8976
rect 3590 8933 3642 8942
rect 3590 8904 3642 8913
rect 3590 8870 3599 8904
rect 3599 8870 3633 8904
rect 3633 8870 3642 8904
rect 3590 8861 3642 8870
rect 4106 9398 4158 9407
rect 4106 9364 4115 9398
rect 4115 9364 4149 9398
rect 4149 9364 4158 9398
rect 4106 9355 4158 9364
rect 4106 9326 4158 9335
rect 4106 9292 4115 9326
rect 4115 9292 4149 9326
rect 4149 9292 4158 9326
rect 4106 9283 4158 9292
rect 4622 9816 4674 9825
rect 4622 9782 4631 9816
rect 4631 9782 4665 9816
rect 4665 9782 4674 9816
rect 4622 9773 4674 9782
rect 4622 9744 4674 9753
rect 4622 9710 4631 9744
rect 4631 9710 4665 9744
rect 4665 9710 4674 9744
rect 4622 9701 4674 9710
rect 4106 8976 4158 8985
rect 4106 8942 4115 8976
rect 4115 8942 4149 8976
rect 4149 8942 4158 8976
rect 4106 8933 4158 8942
rect 4106 8904 4158 8913
rect 4106 8870 4115 8904
rect 4115 8870 4149 8904
rect 4149 8870 4158 8904
rect 4106 8861 4158 8870
rect 4622 9398 4674 9407
rect 4622 9364 4631 9398
rect 4631 9364 4665 9398
rect 4665 9364 4674 9398
rect 4622 9355 4674 9364
rect 4622 9326 4674 9335
rect 4622 9292 4631 9326
rect 4631 9292 4665 9326
rect 4665 9292 4674 9326
rect 4622 9283 4674 9292
rect 4457 9207 4509 9213
rect 4457 9173 4466 9207
rect 4466 9173 4500 9207
rect 4500 9173 4509 9207
rect 4457 9161 4509 9173
rect 4529 9207 4581 9213
rect 4529 9173 4538 9207
rect 4538 9173 4572 9207
rect 4572 9173 4581 9207
rect 4529 9161 4581 9173
rect 4715 9207 4767 9213
rect 4715 9173 4724 9207
rect 4724 9173 4758 9207
rect 4758 9173 4767 9207
rect 4715 9161 4767 9173
rect 4787 9207 4839 9213
rect 4787 9173 4796 9207
rect 4796 9173 4830 9207
rect 4830 9173 4839 9207
rect 4787 9161 4839 9173
rect 4457 9095 4509 9104
rect 4457 9061 4466 9095
rect 4466 9061 4500 9095
rect 4500 9061 4509 9095
rect 4457 9052 4509 9061
rect 4529 9095 4581 9104
rect 4529 9061 4538 9095
rect 4538 9061 4572 9095
rect 4572 9061 4581 9095
rect 4529 9052 4581 9061
rect 4715 9095 4767 9104
rect 4715 9061 4724 9095
rect 4724 9061 4758 9095
rect 4758 9061 4767 9095
rect 4715 9052 4767 9061
rect 4787 9095 4839 9104
rect 4787 9061 4796 9095
rect 4796 9061 4830 9095
rect 4830 9061 4839 9095
rect 4787 9052 4839 9061
rect 3941 8785 3993 8791
rect 3941 8751 3950 8785
rect 3950 8751 3984 8785
rect 3984 8751 3993 8785
rect 3941 8739 3993 8751
rect 4013 8785 4065 8791
rect 4013 8751 4022 8785
rect 4022 8751 4056 8785
rect 4056 8751 4065 8785
rect 4013 8739 4065 8751
rect 4199 8785 4251 8791
rect 4199 8751 4208 8785
rect 4208 8751 4242 8785
rect 4242 8751 4251 8785
rect 4199 8739 4251 8751
rect 4271 8785 4323 8791
rect 4271 8751 4280 8785
rect 4280 8751 4314 8785
rect 4314 8751 4323 8785
rect 4271 8739 4323 8751
rect 4622 8976 4674 8985
rect 4622 8942 4631 8976
rect 4631 8942 4665 8976
rect 4665 8942 4674 8976
rect 4622 8933 4674 8942
rect 4622 8904 4674 8913
rect 4622 8870 4631 8904
rect 4631 8870 4665 8904
rect 4665 8870 4674 8904
rect 4622 8861 4674 8870
rect 2241 8319 2293 8371
rect 3590 8554 3642 8563
rect 3590 8520 3599 8554
rect 3599 8520 3633 8554
rect 3633 8520 3642 8554
rect 3590 8511 3642 8520
rect 3590 8482 3642 8491
rect 3590 8448 3599 8482
rect 3599 8448 3633 8482
rect 3633 8448 3642 8482
rect 3590 8439 3642 8448
rect 3941 8673 3993 8682
rect 3941 8639 3950 8673
rect 3950 8639 3984 8673
rect 3984 8639 3993 8673
rect 3941 8630 3993 8639
rect 4013 8673 4065 8682
rect 4013 8639 4022 8673
rect 4022 8639 4056 8673
rect 4056 8639 4065 8673
rect 4013 8630 4065 8639
rect 4199 8673 4251 8682
rect 4199 8639 4208 8673
rect 4208 8639 4242 8673
rect 4242 8639 4251 8673
rect 4199 8630 4251 8639
rect 4271 8673 4323 8682
rect 4271 8639 4280 8673
rect 4280 8639 4314 8673
rect 4314 8639 4323 8673
rect 4271 8630 4323 8639
rect 3683 8363 3735 8369
rect 3683 8329 3692 8363
rect 3692 8329 3726 8363
rect 3726 8329 3735 8363
rect 3683 8317 3735 8329
rect 3755 8363 3807 8369
rect 3755 8329 3764 8363
rect 3764 8329 3798 8363
rect 3798 8329 3807 8363
rect 3755 8317 3807 8329
rect -834 8022 -782 8031
rect -834 7988 -825 8022
rect -825 7988 -791 8022
rect -791 7988 -782 8022
rect -834 7979 -782 7988
rect -762 8022 -710 8031
rect -762 7988 -753 8022
rect -753 7988 -719 8022
rect -719 7988 -710 8022
rect -762 7979 -710 7988
rect -576 8022 -524 8031
rect -576 7988 -567 8022
rect -567 7988 -533 8022
rect -533 7988 -524 8022
rect -576 7979 -524 7988
rect -504 8022 -452 8031
rect -504 7988 -495 8022
rect -495 7988 -461 8022
rect -461 7988 -452 8022
rect -504 7979 -452 7988
rect -318 8022 -266 8031
rect -318 7988 -309 8022
rect -309 7988 -275 8022
rect -275 7988 -266 8022
rect -318 7979 -266 7988
rect -246 8022 -194 8031
rect -246 7988 -237 8022
rect -237 7988 -203 8022
rect -203 7988 -194 8022
rect -246 7979 -194 7988
rect -60 8022 -8 8031
rect -60 7988 -51 8022
rect -51 7988 -17 8022
rect -17 7988 -8 8022
rect -60 7979 -8 7988
rect 12 8022 64 8031
rect 12 7988 21 8022
rect 21 7988 55 8022
rect 55 7988 64 8022
rect 12 7979 64 7988
rect 198 8022 250 8031
rect 198 7988 207 8022
rect 207 7988 241 8022
rect 241 7988 250 8022
rect 198 7979 250 7988
rect 270 8022 322 8031
rect 270 7988 279 8022
rect 279 7988 313 8022
rect 313 7988 322 8022
rect 270 7979 322 7988
rect 456 8022 508 8031
rect 456 7988 465 8022
rect 465 7988 499 8022
rect 499 7988 508 8022
rect 456 7979 508 7988
rect 528 8022 580 8031
rect 528 7988 537 8022
rect 537 7988 571 8022
rect 571 7988 580 8022
rect 528 7979 580 7988
rect 4106 8554 4158 8563
rect 4106 8520 4115 8554
rect 4115 8520 4149 8554
rect 4149 8520 4158 8554
rect 4106 8511 4158 8520
rect 4106 8482 4158 8491
rect 4106 8448 4115 8482
rect 4115 8448 4149 8482
rect 4149 8448 4158 8482
rect 4106 8439 4158 8448
rect 4622 8554 4674 8563
rect 4622 8520 4631 8554
rect 4631 8520 4665 8554
rect 4665 8520 4674 8554
rect 4622 8511 4674 8520
rect 4622 8482 4674 8491
rect 4622 8448 4631 8482
rect 4631 8448 4665 8482
rect 4665 8448 4674 8482
rect 4622 8439 4674 8448
rect 4457 8363 4509 8369
rect 4457 8329 4466 8363
rect 4466 8329 4500 8363
rect 4500 8329 4509 8363
rect 4457 8317 4509 8329
rect 4529 8363 4581 8369
rect 4529 8329 4538 8363
rect 4538 8329 4572 8363
rect 4572 8329 4581 8363
rect 4529 8317 4581 8329
rect 7351 10551 7403 10560
rect 7351 10517 7360 10551
rect 7360 10517 7394 10551
rect 7394 10517 7403 10551
rect 7351 10508 7403 10517
rect 7423 10551 7475 10560
rect 7423 10517 7432 10551
rect 7432 10517 7466 10551
rect 7466 10517 7475 10551
rect 7423 10508 7475 10517
rect 7351 10443 7403 10452
rect 7351 10409 7360 10443
rect 7360 10409 7394 10443
rect 7394 10409 7403 10443
rect 7351 10400 7403 10409
rect 7423 10443 7475 10452
rect 7423 10409 7432 10443
rect 7432 10409 7466 10443
rect 7466 10409 7475 10443
rect 7423 10400 7475 10409
rect 7609 10551 7661 10560
rect 7609 10517 7618 10551
rect 7618 10517 7652 10551
rect 7652 10517 7661 10551
rect 7609 10508 7661 10517
rect 7681 10551 7733 10560
rect 7681 10517 7690 10551
rect 7690 10517 7724 10551
rect 7724 10517 7733 10551
rect 7681 10508 7733 10517
rect 7609 10443 7661 10452
rect 7609 10409 7618 10443
rect 7618 10409 7652 10443
rect 7652 10409 7661 10443
rect 7609 10400 7661 10409
rect 7681 10443 7733 10452
rect 7681 10409 7690 10443
rect 7690 10409 7724 10443
rect 7724 10409 7733 10443
rect 7681 10400 7733 10409
rect 7351 9679 7403 9688
rect 7351 9645 7360 9679
rect 7360 9645 7394 9679
rect 7394 9645 7403 9679
rect 7351 9636 7403 9645
rect 7423 9679 7475 9688
rect 7423 9645 7432 9679
rect 7432 9645 7466 9679
rect 7466 9645 7475 9679
rect 7423 9636 7475 9645
rect 7351 9571 7403 9580
rect 7351 9537 7360 9571
rect 7360 9537 7394 9571
rect 7394 9537 7403 9571
rect 7351 9528 7403 9537
rect 7423 9571 7475 9580
rect 7423 9537 7432 9571
rect 7432 9537 7466 9571
rect 7466 9537 7475 9571
rect 7423 9528 7475 9537
rect 7867 10551 7919 10560
rect 7867 10517 7876 10551
rect 7876 10517 7910 10551
rect 7910 10517 7919 10551
rect 7867 10508 7919 10517
rect 7939 10551 7991 10560
rect 7939 10517 7948 10551
rect 7948 10517 7982 10551
rect 7982 10517 7991 10551
rect 7939 10508 7991 10517
rect 7867 10443 7919 10452
rect 7867 10409 7876 10443
rect 7876 10409 7910 10443
rect 7910 10409 7919 10443
rect 7867 10400 7919 10409
rect 7939 10443 7991 10452
rect 7939 10409 7948 10443
rect 7948 10409 7982 10443
rect 7982 10409 7991 10443
rect 7939 10400 7991 10409
rect 7609 9679 7661 9688
rect 7609 9645 7618 9679
rect 7618 9645 7652 9679
rect 7652 9645 7661 9679
rect 7609 9636 7661 9645
rect 7681 9679 7733 9688
rect 7681 9645 7690 9679
rect 7690 9645 7724 9679
rect 7724 9645 7733 9679
rect 7681 9636 7733 9645
rect 7609 9571 7661 9580
rect 7609 9537 7618 9571
rect 7618 9537 7652 9571
rect 7652 9537 7661 9571
rect 7609 9528 7661 9537
rect 7681 9571 7733 9580
rect 7681 9537 7690 9571
rect 7690 9537 7724 9571
rect 7724 9537 7733 9571
rect 7681 9528 7733 9537
rect 7351 8807 7403 8816
rect 7351 8773 7360 8807
rect 7360 8773 7394 8807
rect 7394 8773 7403 8807
rect 7351 8764 7403 8773
rect 7423 8807 7475 8816
rect 7423 8773 7432 8807
rect 7432 8773 7466 8807
rect 7466 8773 7475 8807
rect 7423 8764 7475 8773
rect 7351 8699 7403 8708
rect 7351 8665 7360 8699
rect 7360 8665 7394 8699
rect 7394 8665 7403 8699
rect 7351 8656 7403 8665
rect 7423 8699 7475 8708
rect 7423 8665 7432 8699
rect 7432 8665 7466 8699
rect 7466 8665 7475 8699
rect 7423 8656 7475 8665
rect 8125 10551 8177 10560
rect 8125 10517 8134 10551
rect 8134 10517 8168 10551
rect 8168 10517 8177 10551
rect 8125 10508 8177 10517
rect 8197 10551 8249 10560
rect 8197 10517 8206 10551
rect 8206 10517 8240 10551
rect 8240 10517 8249 10551
rect 8197 10508 8249 10517
rect 8125 10443 8177 10452
rect 8125 10409 8134 10443
rect 8134 10409 8168 10443
rect 8168 10409 8177 10443
rect 8125 10400 8177 10409
rect 8197 10443 8249 10452
rect 8197 10409 8206 10443
rect 8206 10409 8240 10443
rect 8240 10409 8249 10443
rect 8197 10400 8249 10409
rect 10024 10777 10076 10829
rect 7867 9679 7919 9688
rect 7867 9645 7876 9679
rect 7876 9645 7910 9679
rect 7910 9645 7919 9679
rect 7867 9636 7919 9645
rect 7939 9679 7991 9688
rect 7939 9645 7948 9679
rect 7948 9645 7982 9679
rect 7982 9645 7991 9679
rect 7939 9636 7991 9645
rect 7867 9571 7919 9580
rect 7867 9537 7876 9571
rect 7876 9537 7910 9571
rect 7910 9537 7919 9571
rect 7867 9528 7919 9537
rect 7939 9571 7991 9580
rect 7939 9537 7948 9571
rect 7948 9537 7982 9571
rect 7982 9537 7991 9571
rect 7939 9528 7991 9537
rect 7609 8807 7661 8816
rect 7609 8773 7618 8807
rect 7618 8773 7652 8807
rect 7652 8773 7661 8807
rect 7609 8764 7661 8773
rect 7681 8807 7733 8816
rect 7681 8773 7690 8807
rect 7690 8773 7724 8807
rect 7724 8773 7733 8807
rect 7681 8764 7733 8773
rect 7609 8699 7661 8708
rect 7609 8665 7618 8699
rect 7618 8665 7652 8699
rect 7652 8665 7661 8699
rect 7609 8656 7661 8665
rect 7681 8699 7733 8708
rect 7681 8665 7690 8699
rect 7690 8665 7724 8699
rect 7724 8665 7733 8699
rect 7681 8656 7733 8665
rect -1350 7604 -1298 7613
rect -1350 7570 -1341 7604
rect -1341 7570 -1307 7604
rect -1307 7570 -1298 7604
rect -1350 7561 -1298 7570
rect -1278 7604 -1226 7613
rect -1278 7570 -1269 7604
rect -1269 7570 -1235 7604
rect -1235 7570 -1226 7604
rect -1278 7561 -1226 7570
rect -1092 7604 -1040 7613
rect -1092 7570 -1083 7604
rect -1083 7570 -1049 7604
rect -1049 7570 -1040 7604
rect -1092 7561 -1040 7570
rect -1020 7604 -968 7613
rect -1020 7570 -1011 7604
rect -1011 7570 -977 7604
rect -977 7570 -968 7604
rect -1020 7561 -968 7570
rect -1185 7485 -1133 7494
rect -1185 7451 -1176 7485
rect -1176 7451 -1142 7485
rect -1142 7451 -1133 7485
rect -1185 7442 -1133 7451
rect -1185 7413 -1133 7422
rect -1185 7379 -1176 7413
rect -1176 7379 -1142 7413
rect -1142 7379 -1133 7413
rect -1185 7370 -1133 7379
rect -669 7903 -617 7912
rect -669 7869 -660 7903
rect -660 7869 -626 7903
rect -626 7869 -617 7903
rect -669 7860 -617 7869
rect -669 7831 -617 7840
rect -669 7797 -660 7831
rect -660 7797 -626 7831
rect -626 7797 -617 7831
rect -669 7788 -617 7797
rect -669 7485 -617 7494
rect -669 7451 -660 7485
rect -660 7451 -626 7485
rect -626 7451 -617 7485
rect -669 7442 -617 7451
rect -669 7413 -617 7422
rect -669 7379 -660 7413
rect -660 7379 -626 7413
rect -626 7379 -617 7413
rect -669 7370 -617 7379
rect -153 7903 -101 7912
rect -153 7869 -144 7903
rect -144 7869 -110 7903
rect -110 7869 -101 7903
rect -153 7860 -101 7869
rect -153 7831 -101 7840
rect -153 7797 -144 7831
rect -144 7797 -110 7831
rect -110 7797 -101 7831
rect -153 7788 -101 7797
rect -318 7604 -266 7613
rect -318 7570 -309 7604
rect -309 7570 -275 7604
rect -275 7570 -266 7604
rect -318 7561 -266 7570
rect -246 7604 -194 7613
rect -246 7570 -237 7604
rect -237 7570 -203 7604
rect -203 7570 -194 7604
rect -246 7561 -194 7570
rect -60 7604 -8 7613
rect -60 7570 -51 7604
rect -51 7570 -17 7604
rect -17 7570 -8 7604
rect -60 7561 -8 7570
rect 12 7604 64 7613
rect 12 7570 21 7604
rect 21 7570 55 7604
rect 55 7570 64 7604
rect 12 7561 64 7570
rect -834 7294 -782 7303
rect -834 7260 -825 7294
rect -825 7260 -791 7294
rect -791 7260 -782 7294
rect -834 7251 -782 7260
rect -762 7294 -710 7303
rect -762 7260 -753 7294
rect -753 7260 -719 7294
rect -719 7260 -710 7294
rect -762 7251 -710 7260
rect -576 7294 -524 7303
rect -576 7260 -567 7294
rect -567 7260 -533 7294
rect -533 7260 -524 7294
rect -576 7251 -524 7260
rect -504 7294 -452 7303
rect -504 7260 -495 7294
rect -495 7260 -461 7294
rect -461 7260 -452 7294
rect -504 7251 -452 7260
rect -153 7485 -101 7494
rect -153 7451 -144 7485
rect -144 7451 -110 7485
rect -110 7451 -101 7485
rect -153 7442 -101 7451
rect -153 7413 -101 7422
rect -153 7379 -144 7413
rect -144 7379 -110 7413
rect -110 7379 -101 7413
rect -153 7370 -101 7379
rect 363 7903 415 7912
rect 363 7869 372 7903
rect 372 7869 406 7903
rect 406 7869 415 7903
rect 363 7860 415 7869
rect 363 7831 415 7840
rect 363 7797 372 7831
rect 372 7797 406 7831
rect 406 7797 415 7831
rect 363 7788 415 7797
rect 363 7485 415 7494
rect 363 7451 372 7485
rect 372 7451 406 7485
rect 406 7451 415 7485
rect 363 7442 415 7451
rect 363 7413 415 7422
rect 363 7379 372 7413
rect 372 7379 406 7413
rect 406 7379 415 7413
rect 363 7370 415 7379
rect 3211 7930 3263 7982
rect 7351 8263 7403 8272
rect 7351 8229 7360 8263
rect 7360 8229 7394 8263
rect 7394 8229 7403 8263
rect 7351 8220 7403 8229
rect 7423 8263 7475 8272
rect 7423 8229 7432 8263
rect 7432 8229 7466 8263
rect 7466 8229 7475 8263
rect 7423 8220 7475 8229
rect 8125 9679 8177 9688
rect 8125 9645 8134 9679
rect 8134 9645 8168 9679
rect 8168 9645 8177 9679
rect 8125 9636 8177 9645
rect 8197 9679 8249 9688
rect 8197 9645 8206 9679
rect 8206 9645 8240 9679
rect 8240 9645 8249 9679
rect 8197 9636 8249 9645
rect 8125 9571 8177 9580
rect 8125 9537 8134 9571
rect 8134 9537 8168 9571
rect 8168 9537 8177 9571
rect 8125 9528 8177 9537
rect 8197 9571 8249 9580
rect 8197 9537 8206 9571
rect 8206 9537 8240 9571
rect 8240 9537 8249 9571
rect 8197 9528 8249 9537
rect 7867 8807 7919 8816
rect 7867 8773 7876 8807
rect 7876 8773 7910 8807
rect 7910 8773 7919 8807
rect 7867 8764 7919 8773
rect 7939 8807 7991 8816
rect 7939 8773 7948 8807
rect 7948 8773 7982 8807
rect 7982 8773 7991 8807
rect 7939 8764 7991 8773
rect 7867 8699 7919 8708
rect 7867 8665 7876 8699
rect 7876 8665 7910 8699
rect 7910 8665 7919 8699
rect 7867 8656 7919 8665
rect 7939 8699 7991 8708
rect 7939 8665 7948 8699
rect 7948 8665 7982 8699
rect 7982 8665 7991 8699
rect 7939 8656 7991 8665
rect 7609 8263 7661 8272
rect 7609 8229 7618 8263
rect 7618 8229 7652 8263
rect 7652 8229 7661 8263
rect 7609 8220 7661 8229
rect 7681 8263 7733 8272
rect 7681 8229 7690 8263
rect 7690 8229 7724 8263
rect 7724 8229 7733 8263
rect 7681 8220 7733 8229
rect 714 7604 766 7613
rect 714 7570 723 7604
rect 723 7570 757 7604
rect 757 7570 766 7604
rect 714 7561 766 7570
rect 786 7604 838 7613
rect 786 7570 795 7604
rect 795 7570 829 7604
rect 829 7570 838 7604
rect 786 7561 838 7570
rect 972 7604 1024 7613
rect 972 7570 981 7604
rect 981 7570 1015 7604
rect 1015 7570 1024 7604
rect 972 7561 1024 7570
rect 1044 7604 1096 7613
rect 1044 7570 1053 7604
rect 1053 7570 1087 7604
rect 1087 7570 1096 7604
rect 1044 7561 1096 7570
rect -1866 7186 -1814 7195
rect -1866 7152 -1857 7186
rect -1857 7152 -1823 7186
rect -1823 7152 -1814 7186
rect -1866 7143 -1814 7152
rect -1794 7186 -1742 7195
rect -1794 7152 -1785 7186
rect -1785 7152 -1751 7186
rect -1751 7152 -1742 7186
rect -1794 7143 -1742 7152
rect -1608 7186 -1556 7195
rect -1608 7152 -1599 7186
rect -1599 7152 -1565 7186
rect -1565 7152 -1556 7186
rect -1608 7143 -1556 7152
rect -1536 7186 -1484 7195
rect -1536 7152 -1527 7186
rect -1527 7152 -1493 7186
rect -1493 7152 -1484 7186
rect -1536 7143 -1484 7152
rect -1701 7067 -1649 7076
rect -1701 7033 -1692 7067
rect -1692 7033 -1658 7067
rect -1658 7033 -1649 7067
rect -1701 7024 -1649 7033
rect -1701 6995 -1649 7004
rect -1701 6961 -1692 6995
rect -1692 6961 -1658 6995
rect -1658 6961 -1649 6995
rect -1701 6952 -1649 6961
rect -1185 7067 -1133 7076
rect -1185 7033 -1176 7067
rect -1176 7033 -1142 7067
rect -1142 7033 -1133 7067
rect -1185 7024 -1133 7033
rect -1185 6995 -1133 7004
rect -1185 6961 -1176 6995
rect -1176 6961 -1142 6995
rect -1142 6961 -1133 6995
rect -1185 6952 -1133 6961
rect 198 7294 250 7303
rect 198 7260 207 7294
rect 207 7260 241 7294
rect 241 7260 250 7294
rect 198 7251 250 7260
rect 270 7294 322 7303
rect 270 7260 279 7294
rect 279 7260 313 7294
rect 313 7260 322 7294
rect 270 7251 322 7260
rect 456 7294 508 7303
rect 456 7260 465 7294
rect 465 7260 499 7294
rect 499 7260 508 7294
rect 456 7251 508 7260
rect 528 7294 580 7303
rect 528 7260 537 7294
rect 537 7260 571 7294
rect 571 7260 580 7294
rect 528 7251 580 7260
rect 879 7485 931 7494
rect 879 7451 888 7485
rect 888 7451 922 7485
rect 922 7451 931 7485
rect 879 7442 931 7451
rect 879 7413 931 7422
rect 879 7379 888 7413
rect 888 7379 922 7413
rect 922 7379 931 7413
rect 879 7370 931 7379
rect 8125 8807 8177 8816
rect 8125 8773 8134 8807
rect 8134 8773 8168 8807
rect 8168 8773 8177 8807
rect 8125 8764 8177 8773
rect 8197 8807 8249 8816
rect 8197 8773 8206 8807
rect 8206 8773 8240 8807
rect 8240 8773 8249 8807
rect 8197 8764 8249 8773
rect 8125 8699 8177 8708
rect 8125 8665 8134 8699
rect 8134 8665 8168 8699
rect 8168 8665 8177 8699
rect 8125 8656 8177 8665
rect 8197 8699 8249 8708
rect 8197 8665 8206 8699
rect 8206 8665 8240 8699
rect 8240 8665 8249 8699
rect 8197 8656 8249 8665
rect 7867 8263 7919 8272
rect 7867 8229 7876 8263
rect 7876 8229 7910 8263
rect 7910 8229 7919 8263
rect 7867 8220 7919 8229
rect 7939 8263 7991 8272
rect 7939 8229 7948 8263
rect 7948 8229 7982 8263
rect 7982 8229 7991 8263
rect 7939 8220 7991 8229
rect 8125 8263 8177 8272
rect 8125 8229 8134 8263
rect 8134 8229 8168 8263
rect 8168 8229 8177 8263
rect 8125 8220 8177 8229
rect 8197 8263 8249 8272
rect 8197 8229 8206 8263
rect 8206 8229 8240 8263
rect 8240 8229 8249 8263
rect 8197 8220 8249 8229
rect -834 7186 -782 7195
rect -834 7152 -825 7186
rect -825 7152 -791 7186
rect -791 7152 -782 7186
rect -834 7143 -782 7152
rect -762 7186 -710 7195
rect -762 7152 -753 7186
rect -753 7152 -719 7186
rect -719 7152 -710 7186
rect -762 7143 -710 7152
rect -576 7186 -524 7195
rect -576 7152 -567 7186
rect -567 7152 -533 7186
rect -533 7152 -524 7186
rect -576 7143 -524 7152
rect -504 7186 -452 7195
rect -504 7152 -495 7186
rect -495 7152 -461 7186
rect -461 7152 -452 7186
rect -504 7143 -452 7152
rect -1350 6876 -1298 6885
rect -1350 6842 -1341 6876
rect -1341 6842 -1307 6876
rect -1307 6842 -1298 6876
rect -1350 6833 -1298 6842
rect -1278 6876 -1226 6885
rect -1278 6842 -1269 6876
rect -1269 6842 -1235 6876
rect -1235 6842 -1226 6876
rect -1278 6833 -1226 6842
rect -1092 6876 -1040 6885
rect -1092 6842 -1083 6876
rect -1083 6842 -1049 6876
rect -1049 6842 -1040 6876
rect -1092 6833 -1040 6842
rect -1020 6876 -968 6885
rect -1020 6842 -1011 6876
rect -1011 6842 -977 6876
rect -977 6842 -968 6876
rect -1020 6833 -968 6842
rect -669 7067 -617 7076
rect -669 7033 -660 7067
rect -660 7033 -626 7067
rect -626 7033 -617 7067
rect -669 7024 -617 7033
rect -669 6995 -617 7004
rect -669 6961 -660 6995
rect -660 6961 -626 6995
rect -626 6961 -617 6995
rect -669 6952 -617 6961
rect -153 7067 -101 7076
rect -153 7033 -144 7067
rect -144 7033 -110 7067
rect -110 7033 -101 7067
rect -153 7024 -101 7033
rect -153 6995 -101 7004
rect -153 6961 -144 6995
rect -144 6961 -110 6995
rect -110 6961 -101 6995
rect -153 6952 -101 6961
rect 198 7186 250 7195
rect 198 7152 207 7186
rect 207 7152 241 7186
rect 241 7152 250 7186
rect 198 7143 250 7152
rect 270 7186 322 7195
rect 270 7152 279 7186
rect 279 7152 313 7186
rect 313 7152 322 7186
rect 270 7143 322 7152
rect 456 7186 508 7195
rect 456 7152 465 7186
rect 465 7152 499 7186
rect 499 7152 508 7186
rect 456 7143 508 7152
rect 528 7186 580 7195
rect 528 7152 537 7186
rect 537 7152 571 7186
rect 571 7152 580 7186
rect 528 7143 580 7152
rect -318 6876 -266 6885
rect -318 6842 -309 6876
rect -309 6842 -275 6876
rect -275 6842 -266 6876
rect -318 6833 -266 6842
rect -246 6876 -194 6885
rect -246 6842 -237 6876
rect -237 6842 -203 6876
rect -203 6842 -194 6876
rect -246 6833 -194 6842
rect -60 6876 -8 6885
rect -60 6842 -51 6876
rect -51 6842 -17 6876
rect -17 6842 -8 6876
rect -60 6833 -8 6842
rect 12 6876 64 6885
rect 12 6842 21 6876
rect 21 6842 55 6876
rect 55 6842 64 6876
rect 12 6833 64 6842
rect -1701 6649 -1649 6658
rect -1701 6615 -1692 6649
rect -1692 6615 -1658 6649
rect -1658 6615 -1649 6649
rect -1701 6606 -1649 6615
rect -1701 6577 -1649 6586
rect -1701 6543 -1692 6577
rect -1692 6543 -1658 6577
rect -1658 6543 -1649 6577
rect -1701 6534 -1649 6543
rect -1350 6768 -1298 6777
rect -1350 6734 -1341 6768
rect -1341 6734 -1307 6768
rect -1307 6734 -1298 6768
rect -1350 6725 -1298 6734
rect -1278 6768 -1226 6777
rect -1278 6734 -1269 6768
rect -1269 6734 -1235 6768
rect -1235 6734 -1226 6768
rect -1278 6725 -1226 6734
rect -1092 6768 -1040 6777
rect -1092 6734 -1083 6768
rect -1083 6734 -1049 6768
rect -1049 6734 -1040 6768
rect -1092 6725 -1040 6734
rect -1020 6768 -968 6777
rect -1020 6734 -1011 6768
rect -1011 6734 -977 6768
rect -977 6734 -968 6768
rect -1020 6725 -968 6734
rect 363 7067 415 7076
rect 363 7033 372 7067
rect 372 7033 406 7067
rect 406 7033 415 7067
rect 363 7024 415 7033
rect 363 6995 415 7004
rect 363 6961 372 6995
rect 372 6961 406 6995
rect 406 6961 415 6995
rect 363 6952 415 6961
rect 879 7067 931 7076
rect 879 7033 888 7067
rect 888 7033 922 7067
rect 922 7033 931 7067
rect 879 7024 931 7033
rect 879 6995 931 7004
rect 879 6961 888 6995
rect 888 6961 922 6995
rect 922 6961 931 6995
rect 879 6952 931 6961
rect 714 6876 766 6885
rect 714 6842 723 6876
rect 723 6842 757 6876
rect 757 6842 766 6876
rect 714 6833 766 6842
rect 786 6876 838 6885
rect 786 6842 795 6876
rect 795 6842 829 6876
rect 829 6842 838 6876
rect 786 6833 838 6842
rect 972 6876 1024 6885
rect 972 6842 981 6876
rect 981 6842 1015 6876
rect 1015 6842 1024 6876
rect 972 6833 1024 6842
rect 1044 6876 1096 6885
rect 1044 6842 1053 6876
rect 1053 6842 1087 6876
rect 1087 6842 1096 6876
rect 1044 6833 1096 6842
rect -1866 6458 -1814 6467
rect -1866 6424 -1857 6458
rect -1857 6424 -1823 6458
rect -1823 6424 -1814 6458
rect -1866 6415 -1814 6424
rect -1794 6458 -1742 6467
rect -1794 6424 -1785 6458
rect -1785 6424 -1751 6458
rect -1751 6424 -1742 6458
rect -1794 6415 -1742 6424
rect -1608 6458 -1556 6467
rect -1608 6424 -1599 6458
rect -1599 6424 -1565 6458
rect -1565 6424 -1556 6458
rect -1608 6415 -1556 6424
rect -1536 6458 -1484 6467
rect -1536 6424 -1527 6458
rect -1527 6424 -1493 6458
rect -1493 6424 -1484 6458
rect -1536 6415 -1484 6424
rect -1866 6350 -1814 6359
rect -1866 6316 -1857 6350
rect -1857 6316 -1823 6350
rect -1823 6316 -1814 6350
rect -1866 6307 -1814 6316
rect -1794 6350 -1742 6359
rect -1794 6316 -1785 6350
rect -1785 6316 -1751 6350
rect -1751 6316 -1742 6350
rect -1794 6307 -1742 6316
rect -1608 6350 -1556 6359
rect -1608 6316 -1599 6350
rect -1599 6316 -1565 6350
rect -1565 6316 -1556 6350
rect -1608 6307 -1556 6316
rect -1536 6350 -1484 6359
rect -1536 6316 -1527 6350
rect -1527 6316 -1493 6350
rect -1493 6316 -1484 6350
rect -1536 6307 -1484 6316
rect -1701 6231 -1649 6240
rect -1701 6197 -1692 6231
rect -1692 6197 -1658 6231
rect -1658 6197 -1649 6231
rect -1701 6188 -1649 6197
rect -1701 6159 -1649 6168
rect -1701 6125 -1692 6159
rect -1692 6125 -1658 6159
rect -1658 6125 -1649 6159
rect -1701 6116 -1649 6125
rect -1185 6649 -1133 6658
rect -1185 6615 -1176 6649
rect -1176 6615 -1142 6649
rect -1142 6615 -1133 6649
rect -1185 6606 -1133 6615
rect -1185 6577 -1133 6586
rect -1185 6543 -1176 6577
rect -1176 6543 -1142 6577
rect -1142 6543 -1133 6577
rect -1185 6534 -1133 6543
rect -1701 5813 -1649 5822
rect -1701 5779 -1692 5813
rect -1692 5779 -1658 5813
rect -1658 5779 -1649 5813
rect -1701 5770 -1649 5779
rect -1701 5741 -1649 5750
rect -1701 5707 -1692 5741
rect -1692 5707 -1658 5741
rect -1658 5707 -1649 5741
rect -1701 5698 -1649 5707
rect -1185 6231 -1133 6240
rect -1185 6197 -1176 6231
rect -1176 6197 -1142 6231
rect -1142 6197 -1133 6231
rect -1185 6188 -1133 6197
rect -1185 6159 -1133 6168
rect -1185 6125 -1176 6159
rect -1176 6125 -1142 6159
rect -1142 6125 -1133 6159
rect -1185 6116 -1133 6125
rect -669 6649 -617 6658
rect -669 6615 -660 6649
rect -660 6615 -626 6649
rect -626 6615 -617 6649
rect -669 6606 -617 6615
rect -669 6577 -617 6586
rect -669 6543 -660 6577
rect -660 6543 -626 6577
rect -626 6543 -617 6577
rect -669 6534 -617 6543
rect -318 6768 -266 6777
rect -318 6734 -309 6768
rect -309 6734 -275 6768
rect -275 6734 -266 6768
rect -318 6725 -266 6734
rect -246 6768 -194 6777
rect -246 6734 -237 6768
rect -237 6734 -203 6768
rect -203 6734 -194 6768
rect -246 6725 -194 6734
rect -60 6768 -8 6777
rect -60 6734 -51 6768
rect -51 6734 -17 6768
rect -17 6734 -8 6768
rect -60 6725 -8 6734
rect 12 6768 64 6777
rect 12 6734 21 6768
rect 21 6734 55 6768
rect 55 6734 64 6768
rect 12 6725 64 6734
rect -834 6458 -782 6467
rect -834 6424 -825 6458
rect -825 6424 -791 6458
rect -791 6424 -782 6458
rect -834 6415 -782 6424
rect -762 6458 -710 6467
rect -762 6424 -753 6458
rect -753 6424 -719 6458
rect -719 6424 -710 6458
rect -762 6415 -710 6424
rect -576 6458 -524 6467
rect -576 6424 -567 6458
rect -567 6424 -533 6458
rect -533 6424 -524 6458
rect -576 6415 -524 6424
rect -504 6458 -452 6467
rect -504 6424 -495 6458
rect -495 6424 -461 6458
rect -461 6424 -452 6458
rect -504 6415 -452 6424
rect -834 6350 -782 6359
rect -834 6316 -825 6350
rect -825 6316 -791 6350
rect -791 6316 -782 6350
rect -834 6307 -782 6316
rect -762 6350 -710 6359
rect -762 6316 -753 6350
rect -753 6316 -719 6350
rect -719 6316 -710 6350
rect -762 6307 -710 6316
rect -576 6350 -524 6359
rect -576 6316 -567 6350
rect -567 6316 -533 6350
rect -533 6316 -524 6350
rect -576 6307 -524 6316
rect -504 6350 -452 6359
rect -504 6316 -495 6350
rect -495 6316 -461 6350
rect -461 6316 -452 6350
rect -504 6307 -452 6316
rect -1350 6040 -1298 6049
rect -1350 6006 -1341 6040
rect -1341 6006 -1307 6040
rect -1307 6006 -1298 6040
rect -1350 5997 -1298 6006
rect -1278 6040 -1226 6049
rect -1278 6006 -1269 6040
rect -1269 6006 -1235 6040
rect -1235 6006 -1226 6040
rect -1278 5997 -1226 6006
rect -1092 6040 -1040 6049
rect -1092 6006 -1083 6040
rect -1083 6006 -1049 6040
rect -1049 6006 -1040 6040
rect -1092 5997 -1040 6006
rect -1020 6040 -968 6049
rect -1020 6006 -1011 6040
rect -1011 6006 -977 6040
rect -977 6006 -968 6040
rect -1020 5997 -968 6006
rect -1350 5932 -1298 5941
rect -1350 5898 -1341 5932
rect -1341 5898 -1307 5932
rect -1307 5898 -1298 5932
rect -1350 5889 -1298 5898
rect -1278 5932 -1226 5941
rect -1278 5898 -1269 5932
rect -1269 5898 -1235 5932
rect -1235 5898 -1226 5932
rect -1278 5889 -1226 5898
rect -1092 5932 -1040 5941
rect -1092 5898 -1083 5932
rect -1083 5898 -1049 5932
rect -1049 5898 -1040 5932
rect -1092 5889 -1040 5898
rect -1020 5932 -968 5941
rect -1020 5898 -1011 5932
rect -1011 5898 -977 5932
rect -977 5898 -968 5932
rect -1020 5889 -968 5898
rect -1866 5622 -1814 5631
rect -1866 5588 -1857 5622
rect -1857 5588 -1823 5622
rect -1823 5588 -1814 5622
rect -1866 5579 -1814 5588
rect -1794 5622 -1742 5631
rect -1794 5588 -1785 5622
rect -1785 5588 -1751 5622
rect -1751 5588 -1742 5622
rect -1794 5579 -1742 5588
rect -1608 5622 -1556 5631
rect -1608 5588 -1599 5622
rect -1599 5588 -1565 5622
rect -1565 5588 -1556 5622
rect -1608 5579 -1556 5588
rect -1536 5622 -1484 5631
rect -1536 5588 -1527 5622
rect -1527 5588 -1493 5622
rect -1493 5588 -1484 5622
rect -1536 5579 -1484 5588
rect -1866 5514 -1814 5523
rect -1866 5480 -1857 5514
rect -1857 5480 -1823 5514
rect -1823 5480 -1814 5514
rect -1866 5471 -1814 5480
rect -1794 5514 -1742 5523
rect -1794 5480 -1785 5514
rect -1785 5480 -1751 5514
rect -1751 5480 -1742 5514
rect -1794 5471 -1742 5480
rect -1608 5514 -1556 5523
rect -1608 5480 -1599 5514
rect -1599 5480 -1565 5514
rect -1565 5480 -1556 5514
rect -1608 5471 -1556 5480
rect -1536 5514 -1484 5523
rect -1536 5480 -1527 5514
rect -1527 5480 -1493 5514
rect -1493 5480 -1484 5514
rect -1536 5471 -1484 5480
rect -1701 5395 -1649 5404
rect -1701 5361 -1692 5395
rect -1692 5361 -1658 5395
rect -1658 5361 -1649 5395
rect -1701 5352 -1649 5361
rect -1701 5323 -1649 5332
rect -1701 5289 -1692 5323
rect -1692 5289 -1658 5323
rect -1658 5289 -1649 5323
rect -1701 5280 -1649 5289
rect -1185 5813 -1133 5822
rect -1185 5779 -1176 5813
rect -1176 5779 -1142 5813
rect -1142 5779 -1133 5813
rect -1185 5770 -1133 5779
rect -1185 5741 -1133 5750
rect -1185 5707 -1176 5741
rect -1176 5707 -1142 5741
rect -1142 5707 -1133 5741
rect -1185 5698 -1133 5707
rect -669 6231 -617 6240
rect -669 6197 -660 6231
rect -660 6197 -626 6231
rect -626 6197 -617 6231
rect -669 6188 -617 6197
rect -669 6159 -617 6168
rect -669 6125 -660 6159
rect -660 6125 -626 6159
rect -626 6125 -617 6159
rect -669 6116 -617 6125
rect -153 6649 -101 6658
rect -153 6615 -144 6649
rect -144 6615 -110 6649
rect -110 6615 -101 6649
rect -153 6606 -101 6615
rect -153 6577 -101 6586
rect -153 6543 -144 6577
rect -144 6543 -110 6577
rect -110 6543 -101 6577
rect -153 6534 -101 6543
rect -1701 4977 -1649 4986
rect -1701 4943 -1692 4977
rect -1692 4943 -1658 4977
rect -1658 4943 -1649 4977
rect -1701 4934 -1649 4943
rect -1701 4905 -1649 4914
rect -1701 4871 -1692 4905
rect -1692 4871 -1658 4905
rect -1658 4871 -1649 4905
rect -1701 4862 -1649 4871
rect -1185 5395 -1133 5404
rect -1185 5361 -1176 5395
rect -1176 5361 -1142 5395
rect -1142 5361 -1133 5395
rect -1185 5352 -1133 5361
rect -1185 5323 -1133 5332
rect -1185 5289 -1176 5323
rect -1176 5289 -1142 5323
rect -1142 5289 -1133 5323
rect -1185 5280 -1133 5289
rect -669 5813 -617 5822
rect -669 5779 -660 5813
rect -660 5779 -626 5813
rect -626 5779 -617 5813
rect -669 5770 -617 5779
rect -669 5741 -617 5750
rect -669 5707 -660 5741
rect -660 5707 -626 5741
rect -626 5707 -617 5741
rect -669 5698 -617 5707
rect -153 6231 -101 6240
rect -153 6197 -144 6231
rect -144 6197 -110 6231
rect -110 6197 -101 6231
rect -153 6188 -101 6197
rect -153 6159 -101 6168
rect -153 6125 -144 6159
rect -144 6125 -110 6159
rect -110 6125 -101 6159
rect -153 6116 -101 6125
rect 363 6649 415 6658
rect 363 6615 372 6649
rect 372 6615 406 6649
rect 406 6615 415 6649
rect 363 6606 415 6615
rect 363 6577 415 6586
rect 363 6543 372 6577
rect 372 6543 406 6577
rect 406 6543 415 6577
rect 363 6534 415 6543
rect 714 6768 766 6777
rect 714 6734 723 6768
rect 723 6734 757 6768
rect 757 6734 766 6768
rect 714 6725 766 6734
rect 786 6768 838 6777
rect 786 6734 795 6768
rect 795 6734 829 6768
rect 829 6734 838 6768
rect 786 6725 838 6734
rect 972 6768 1024 6777
rect 972 6734 981 6768
rect 981 6734 1015 6768
rect 1015 6734 1024 6768
rect 972 6725 1024 6734
rect 1044 6768 1096 6777
rect 1044 6734 1053 6768
rect 1053 6734 1087 6768
rect 1087 6734 1096 6768
rect 1044 6725 1096 6734
rect 198 6458 250 6467
rect 198 6424 207 6458
rect 207 6424 241 6458
rect 241 6424 250 6458
rect 198 6415 250 6424
rect 270 6458 322 6467
rect 270 6424 279 6458
rect 279 6424 313 6458
rect 313 6424 322 6458
rect 270 6415 322 6424
rect 456 6458 508 6467
rect 456 6424 465 6458
rect 465 6424 499 6458
rect 499 6424 508 6458
rect 456 6415 508 6424
rect 528 6458 580 6467
rect 528 6424 537 6458
rect 537 6424 571 6458
rect 571 6424 580 6458
rect 528 6415 580 6424
rect 198 6350 250 6359
rect 198 6316 207 6350
rect 207 6316 241 6350
rect 241 6316 250 6350
rect 198 6307 250 6316
rect 270 6350 322 6359
rect 270 6316 279 6350
rect 279 6316 313 6350
rect 313 6316 322 6350
rect 270 6307 322 6316
rect 456 6350 508 6359
rect 456 6316 465 6350
rect 465 6316 499 6350
rect 499 6316 508 6350
rect 456 6307 508 6316
rect 528 6350 580 6359
rect 528 6316 537 6350
rect 537 6316 571 6350
rect 571 6316 580 6350
rect 528 6307 580 6316
rect -318 6040 -266 6049
rect -318 6006 -309 6040
rect -309 6006 -275 6040
rect -275 6006 -266 6040
rect -318 5997 -266 6006
rect -246 6040 -194 6049
rect -246 6006 -237 6040
rect -237 6006 -203 6040
rect -203 6006 -194 6040
rect -246 5997 -194 6006
rect -60 6040 -8 6049
rect -60 6006 -51 6040
rect -51 6006 -17 6040
rect -17 6006 -8 6040
rect -60 5997 -8 6006
rect 12 6040 64 6049
rect 12 6006 21 6040
rect 21 6006 55 6040
rect 55 6006 64 6040
rect 12 5997 64 6006
rect -318 5932 -266 5941
rect -318 5898 -309 5932
rect -309 5898 -275 5932
rect -275 5898 -266 5932
rect -318 5889 -266 5898
rect -246 5932 -194 5941
rect -246 5898 -237 5932
rect -237 5898 -203 5932
rect -203 5898 -194 5932
rect -246 5889 -194 5898
rect -60 5932 -8 5941
rect -60 5898 -51 5932
rect -51 5898 -17 5932
rect -17 5898 -8 5932
rect -60 5889 -8 5898
rect 12 5932 64 5941
rect 12 5898 21 5932
rect 21 5898 55 5932
rect 55 5898 64 5932
rect 12 5889 64 5898
rect -834 5622 -782 5631
rect -834 5588 -825 5622
rect -825 5588 -791 5622
rect -791 5588 -782 5622
rect -834 5579 -782 5588
rect -762 5622 -710 5631
rect -762 5588 -753 5622
rect -753 5588 -719 5622
rect -719 5588 -710 5622
rect -762 5579 -710 5588
rect -576 5622 -524 5631
rect -576 5588 -567 5622
rect -567 5588 -533 5622
rect -533 5588 -524 5622
rect -576 5579 -524 5588
rect -504 5622 -452 5631
rect -504 5588 -495 5622
rect -495 5588 -461 5622
rect -461 5588 -452 5622
rect -504 5579 -452 5588
rect -834 5514 -782 5523
rect -834 5480 -825 5514
rect -825 5480 -791 5514
rect -791 5480 -782 5514
rect -834 5471 -782 5480
rect -762 5514 -710 5523
rect -762 5480 -753 5514
rect -753 5480 -719 5514
rect -719 5480 -710 5514
rect -762 5471 -710 5480
rect -576 5514 -524 5523
rect -576 5480 -567 5514
rect -567 5480 -533 5514
rect -533 5480 -524 5514
rect -576 5471 -524 5480
rect -504 5514 -452 5523
rect -504 5480 -495 5514
rect -495 5480 -461 5514
rect -461 5480 -452 5514
rect -504 5471 -452 5480
rect -1350 5204 -1298 5213
rect -1350 5170 -1341 5204
rect -1341 5170 -1307 5204
rect -1307 5170 -1298 5204
rect -1350 5161 -1298 5170
rect -1278 5204 -1226 5213
rect -1278 5170 -1269 5204
rect -1269 5170 -1235 5204
rect -1235 5170 -1226 5204
rect -1278 5161 -1226 5170
rect -1092 5204 -1040 5213
rect -1092 5170 -1083 5204
rect -1083 5170 -1049 5204
rect -1049 5170 -1040 5204
rect -1092 5161 -1040 5170
rect -1020 5204 -968 5213
rect -1020 5170 -1011 5204
rect -1011 5170 -977 5204
rect -977 5170 -968 5204
rect -1020 5161 -968 5170
rect -1350 5096 -1298 5105
rect -1350 5062 -1341 5096
rect -1341 5062 -1307 5096
rect -1307 5062 -1298 5096
rect -1350 5053 -1298 5062
rect -1278 5096 -1226 5105
rect -1278 5062 -1269 5096
rect -1269 5062 -1235 5096
rect -1235 5062 -1226 5096
rect -1278 5053 -1226 5062
rect -1092 5096 -1040 5105
rect -1092 5062 -1083 5096
rect -1083 5062 -1049 5096
rect -1049 5062 -1040 5096
rect -1092 5053 -1040 5062
rect -1020 5096 -968 5105
rect -1020 5062 -1011 5096
rect -1011 5062 -977 5096
rect -977 5062 -968 5096
rect -1020 5053 -968 5062
rect -1866 4786 -1814 4795
rect -1866 4752 -1857 4786
rect -1857 4752 -1823 4786
rect -1823 4752 -1814 4786
rect -1866 4743 -1814 4752
rect -1794 4786 -1742 4795
rect -1794 4752 -1785 4786
rect -1785 4752 -1751 4786
rect -1751 4752 -1742 4786
rect -1794 4743 -1742 4752
rect -1608 4786 -1556 4795
rect -1608 4752 -1599 4786
rect -1599 4752 -1565 4786
rect -1565 4752 -1556 4786
rect -1608 4743 -1556 4752
rect -1536 4786 -1484 4795
rect -1536 4752 -1527 4786
rect -1527 4752 -1493 4786
rect -1493 4752 -1484 4786
rect -1536 4743 -1484 4752
rect -1866 4678 -1814 4687
rect -1866 4644 -1857 4678
rect -1857 4644 -1823 4678
rect -1823 4644 -1814 4678
rect -1866 4635 -1814 4644
rect -1794 4678 -1742 4687
rect -1794 4644 -1785 4678
rect -1785 4644 -1751 4678
rect -1751 4644 -1742 4678
rect -1794 4635 -1742 4644
rect -1608 4678 -1556 4687
rect -1608 4644 -1599 4678
rect -1599 4644 -1565 4678
rect -1565 4644 -1556 4678
rect -1608 4635 -1556 4644
rect -1536 4678 -1484 4687
rect -1536 4644 -1527 4678
rect -1527 4644 -1493 4678
rect -1493 4644 -1484 4678
rect -1536 4635 -1484 4644
rect -1701 4559 -1649 4568
rect -1701 4525 -1692 4559
rect -1692 4525 -1658 4559
rect -1658 4525 -1649 4559
rect -1701 4516 -1649 4525
rect -1701 4487 -1649 4496
rect -1701 4453 -1692 4487
rect -1692 4453 -1658 4487
rect -1658 4453 -1649 4487
rect -1701 4444 -1649 4453
rect -1185 4977 -1133 4986
rect -1185 4943 -1176 4977
rect -1176 4943 -1142 4977
rect -1142 4943 -1133 4977
rect -1185 4934 -1133 4943
rect -1185 4905 -1133 4914
rect -1185 4871 -1176 4905
rect -1176 4871 -1142 4905
rect -1142 4871 -1133 4905
rect -1185 4862 -1133 4871
rect -669 5395 -617 5404
rect -669 5361 -660 5395
rect -660 5361 -626 5395
rect -626 5361 -617 5395
rect -669 5352 -617 5361
rect -669 5323 -617 5332
rect -669 5289 -660 5323
rect -660 5289 -626 5323
rect -626 5289 -617 5323
rect -669 5280 -617 5289
rect -153 5813 -101 5822
rect -153 5779 -144 5813
rect -144 5779 -110 5813
rect -110 5779 -101 5813
rect -153 5770 -101 5779
rect -153 5741 -101 5750
rect -153 5707 -144 5741
rect -144 5707 -110 5741
rect -110 5707 -101 5741
rect -153 5698 -101 5707
rect 363 6231 415 6240
rect 363 6197 372 6231
rect 372 6197 406 6231
rect 406 6197 415 6231
rect 363 6188 415 6197
rect 363 6159 415 6168
rect 363 6125 372 6159
rect 372 6125 406 6159
rect 406 6125 415 6159
rect 363 6116 415 6125
rect 879 6649 931 6658
rect 879 6615 888 6649
rect 888 6615 922 6649
rect 922 6615 931 6649
rect 879 6606 931 6615
rect 879 6577 931 6586
rect 879 6543 888 6577
rect 888 6543 922 6577
rect 922 6543 931 6577
rect 879 6534 931 6543
rect -1185 4559 -1133 4568
rect -1185 4525 -1176 4559
rect -1176 4525 -1142 4559
rect -1142 4525 -1133 4559
rect -1185 4516 -1133 4525
rect -1185 4487 -1133 4496
rect -1185 4453 -1176 4487
rect -1176 4453 -1142 4487
rect -1142 4453 -1133 4487
rect -1185 4444 -1133 4453
rect -669 4977 -617 4986
rect -669 4943 -660 4977
rect -660 4943 -626 4977
rect -626 4943 -617 4977
rect -669 4934 -617 4943
rect -669 4905 -617 4914
rect -669 4871 -660 4905
rect -660 4871 -626 4905
rect -626 4871 -617 4905
rect -669 4862 -617 4871
rect -153 5395 -101 5404
rect -153 5361 -144 5395
rect -144 5361 -110 5395
rect -110 5361 -101 5395
rect -153 5352 -101 5361
rect -153 5323 -101 5332
rect -153 5289 -144 5323
rect -144 5289 -110 5323
rect -110 5289 -101 5323
rect -153 5280 -101 5289
rect 363 5813 415 5822
rect 363 5779 372 5813
rect 372 5779 406 5813
rect 406 5779 415 5813
rect 363 5770 415 5779
rect 363 5741 415 5750
rect 363 5707 372 5741
rect 372 5707 406 5741
rect 406 5707 415 5741
rect 363 5698 415 5707
rect 879 6231 931 6240
rect 879 6197 888 6231
rect 888 6197 922 6231
rect 922 6197 931 6231
rect 879 6188 931 6197
rect 879 6159 931 6168
rect 879 6125 888 6159
rect 888 6125 922 6159
rect 922 6125 931 6159
rect 879 6116 931 6125
rect 714 6040 766 6049
rect 714 6006 723 6040
rect 723 6006 757 6040
rect 757 6006 766 6040
rect 714 5997 766 6006
rect 786 6040 838 6049
rect 786 6006 795 6040
rect 795 6006 829 6040
rect 829 6006 838 6040
rect 786 5997 838 6006
rect 972 6040 1024 6049
rect 972 6006 981 6040
rect 981 6006 1015 6040
rect 1015 6006 1024 6040
rect 972 5997 1024 6006
rect 1044 6040 1096 6049
rect 1044 6006 1053 6040
rect 1053 6006 1087 6040
rect 1087 6006 1096 6040
rect 1044 5997 1096 6006
rect 714 5932 766 5941
rect 714 5898 723 5932
rect 723 5898 757 5932
rect 757 5898 766 5932
rect 714 5889 766 5898
rect 786 5932 838 5941
rect 786 5898 795 5932
rect 795 5898 829 5932
rect 829 5898 838 5932
rect 786 5889 838 5898
rect 972 5932 1024 5941
rect 972 5898 981 5932
rect 981 5898 1015 5932
rect 1015 5898 1024 5932
rect 972 5889 1024 5898
rect 1044 5932 1096 5941
rect 1044 5898 1053 5932
rect 1053 5898 1087 5932
rect 1087 5898 1096 5932
rect 1044 5889 1096 5898
rect 198 5622 250 5631
rect 198 5588 207 5622
rect 207 5588 241 5622
rect 241 5588 250 5622
rect 198 5579 250 5588
rect 270 5622 322 5631
rect 270 5588 279 5622
rect 279 5588 313 5622
rect 313 5588 322 5622
rect 270 5579 322 5588
rect 456 5622 508 5631
rect 456 5588 465 5622
rect 465 5588 499 5622
rect 499 5588 508 5622
rect 456 5579 508 5588
rect 528 5622 580 5631
rect 528 5588 537 5622
rect 537 5588 571 5622
rect 571 5588 580 5622
rect 528 5579 580 5588
rect 198 5514 250 5523
rect 198 5480 207 5514
rect 207 5480 241 5514
rect 241 5480 250 5514
rect 198 5471 250 5480
rect 270 5514 322 5523
rect 270 5480 279 5514
rect 279 5480 313 5514
rect 313 5480 322 5514
rect 270 5471 322 5480
rect 456 5514 508 5523
rect 456 5480 465 5514
rect 465 5480 499 5514
rect 499 5480 508 5514
rect 456 5471 508 5480
rect 528 5514 580 5523
rect 528 5480 537 5514
rect 537 5480 571 5514
rect 571 5480 580 5514
rect 528 5471 580 5480
rect -318 5204 -266 5213
rect -318 5170 -309 5204
rect -309 5170 -275 5204
rect -275 5170 -266 5204
rect -318 5161 -266 5170
rect -246 5204 -194 5213
rect -246 5170 -237 5204
rect -237 5170 -203 5204
rect -203 5170 -194 5204
rect -246 5161 -194 5170
rect -60 5204 -8 5213
rect -60 5170 -51 5204
rect -51 5170 -17 5204
rect -17 5170 -8 5204
rect -60 5161 -8 5170
rect 12 5204 64 5213
rect 12 5170 21 5204
rect 21 5170 55 5204
rect 55 5170 64 5204
rect 12 5161 64 5170
rect -318 5096 -266 5105
rect -318 5062 -309 5096
rect -309 5062 -275 5096
rect -275 5062 -266 5096
rect -318 5053 -266 5062
rect -246 5096 -194 5105
rect -246 5062 -237 5096
rect -237 5062 -203 5096
rect -203 5062 -194 5096
rect -246 5053 -194 5062
rect -60 5096 -8 5105
rect -60 5062 -51 5096
rect -51 5062 -17 5096
rect -17 5062 -8 5096
rect -60 5053 -8 5062
rect 12 5096 64 5105
rect 12 5062 21 5096
rect 21 5062 55 5096
rect 55 5062 64 5096
rect 12 5053 64 5062
rect -834 4786 -782 4795
rect -834 4752 -825 4786
rect -825 4752 -791 4786
rect -791 4752 -782 4786
rect -834 4743 -782 4752
rect -762 4786 -710 4795
rect -762 4752 -753 4786
rect -753 4752 -719 4786
rect -719 4752 -710 4786
rect -762 4743 -710 4752
rect -576 4786 -524 4795
rect -576 4752 -567 4786
rect -567 4752 -533 4786
rect -533 4752 -524 4786
rect -576 4743 -524 4752
rect -504 4786 -452 4795
rect -504 4752 -495 4786
rect -495 4752 -461 4786
rect -461 4752 -452 4786
rect -504 4743 -452 4752
rect -834 4678 -782 4687
rect -834 4644 -825 4678
rect -825 4644 -791 4678
rect -791 4644 -782 4678
rect -834 4635 -782 4644
rect -762 4678 -710 4687
rect -762 4644 -753 4678
rect -753 4644 -719 4678
rect -719 4644 -710 4678
rect -762 4635 -710 4644
rect -576 4678 -524 4687
rect -576 4644 -567 4678
rect -567 4644 -533 4678
rect -533 4644 -524 4678
rect -576 4635 -524 4644
rect -504 4678 -452 4687
rect -504 4644 -495 4678
rect -495 4644 -461 4678
rect -461 4644 -452 4678
rect -504 4635 -452 4644
rect -1350 4368 -1298 4377
rect -1350 4334 -1341 4368
rect -1341 4334 -1307 4368
rect -1307 4334 -1298 4368
rect -1350 4325 -1298 4334
rect -1278 4368 -1226 4377
rect -1278 4334 -1269 4368
rect -1269 4334 -1235 4368
rect -1235 4334 -1226 4368
rect -1278 4325 -1226 4334
rect -1092 4368 -1040 4377
rect -1092 4334 -1083 4368
rect -1083 4334 -1049 4368
rect -1049 4334 -1040 4368
rect -1092 4325 -1040 4334
rect -1020 4368 -968 4377
rect -1020 4334 -1011 4368
rect -1011 4334 -977 4368
rect -977 4334 -968 4368
rect -1020 4325 -968 4334
rect -1350 4260 -1298 4269
rect -1350 4226 -1341 4260
rect -1341 4226 -1307 4260
rect -1307 4226 -1298 4260
rect -1350 4217 -1298 4226
rect -1278 4260 -1226 4269
rect -1278 4226 -1269 4260
rect -1269 4226 -1235 4260
rect -1235 4226 -1226 4260
rect -1278 4217 -1226 4226
rect -1092 4260 -1040 4269
rect -1092 4226 -1083 4260
rect -1083 4226 -1049 4260
rect -1049 4226 -1040 4260
rect -1092 4217 -1040 4226
rect -1020 4260 -968 4269
rect -1020 4226 -1011 4260
rect -1011 4226 -977 4260
rect -977 4226 -968 4260
rect -1020 4217 -968 4226
rect -1185 4141 -1133 4150
rect -1185 4107 -1176 4141
rect -1176 4107 -1142 4141
rect -1142 4107 -1133 4141
rect -1185 4098 -1133 4107
rect -1185 4069 -1133 4078
rect -1185 4035 -1176 4069
rect -1176 4035 -1142 4069
rect -1142 4035 -1133 4069
rect -1185 4026 -1133 4035
rect -669 4559 -617 4568
rect -669 4525 -660 4559
rect -660 4525 -626 4559
rect -626 4525 -617 4559
rect -669 4516 -617 4525
rect -669 4487 -617 4496
rect -669 4453 -660 4487
rect -660 4453 -626 4487
rect -626 4453 -617 4487
rect -669 4444 -617 4453
rect -153 4977 -101 4986
rect -153 4943 -144 4977
rect -144 4943 -110 4977
rect -110 4943 -101 4977
rect -153 4934 -101 4943
rect -153 4905 -101 4914
rect -153 4871 -144 4905
rect -144 4871 -110 4905
rect -110 4871 -101 4905
rect -153 4862 -101 4871
rect 363 5395 415 5404
rect 363 5361 372 5395
rect 372 5361 406 5395
rect 406 5361 415 5395
rect 363 5352 415 5361
rect 363 5323 415 5332
rect 363 5289 372 5323
rect 372 5289 406 5323
rect 406 5289 415 5323
rect 363 5280 415 5289
rect 879 5813 931 5822
rect 879 5779 888 5813
rect 888 5779 922 5813
rect 922 5779 931 5813
rect 879 5770 931 5779
rect 879 5741 931 5750
rect 879 5707 888 5741
rect 888 5707 922 5741
rect 922 5707 931 5741
rect 879 5698 931 5707
rect -834 4260 -782 4269
rect -834 4226 -825 4260
rect -825 4226 -791 4260
rect -791 4226 -782 4260
rect -834 4217 -782 4226
rect -762 4260 -710 4269
rect -762 4226 -753 4260
rect -753 4226 -719 4260
rect -719 4226 -710 4260
rect -762 4217 -710 4226
rect -576 4260 -524 4269
rect -576 4226 -567 4260
rect -567 4226 -533 4260
rect -533 4226 -524 4260
rect -576 4217 -524 4226
rect -504 4260 -452 4269
rect -504 4226 -495 4260
rect -495 4226 -461 4260
rect -461 4226 -452 4260
rect -504 4217 -452 4226
rect -669 4141 -617 4150
rect -669 4107 -660 4141
rect -660 4107 -626 4141
rect -626 4107 -617 4141
rect -669 4098 -617 4107
rect -669 4069 -617 4078
rect -669 4035 -660 4069
rect -660 4035 -626 4069
rect -626 4035 -617 4069
rect -669 4026 -617 4035
rect -153 4559 -101 4568
rect -153 4525 -144 4559
rect -144 4525 -110 4559
rect -110 4525 -101 4559
rect -153 4516 -101 4525
rect -153 4487 -101 4496
rect -153 4453 -144 4487
rect -144 4453 -110 4487
rect -110 4453 -101 4487
rect -153 4444 -101 4453
rect 363 4977 415 4986
rect 363 4943 372 4977
rect 372 4943 406 4977
rect 406 4943 415 4977
rect 363 4934 415 4943
rect 363 4905 415 4914
rect 363 4871 372 4905
rect 372 4871 406 4905
rect 406 4871 415 4905
rect 363 4862 415 4871
rect 879 5395 931 5404
rect 879 5361 888 5395
rect 888 5361 922 5395
rect 922 5361 931 5395
rect 879 5352 931 5361
rect 879 5323 931 5332
rect 879 5289 888 5323
rect 888 5289 922 5323
rect 922 5289 931 5323
rect 879 5280 931 5289
rect 714 5204 766 5213
rect 714 5170 723 5204
rect 723 5170 757 5204
rect 757 5170 766 5204
rect 714 5161 766 5170
rect 786 5204 838 5213
rect 786 5170 795 5204
rect 795 5170 829 5204
rect 829 5170 838 5204
rect 786 5161 838 5170
rect 972 5204 1024 5213
rect 972 5170 981 5204
rect 981 5170 1015 5204
rect 1015 5170 1024 5204
rect 972 5161 1024 5170
rect 1044 5204 1096 5213
rect 1044 5170 1053 5204
rect 1053 5170 1087 5204
rect 1087 5170 1096 5204
rect 1044 5161 1096 5170
rect 714 5096 766 5105
rect 714 5062 723 5096
rect 723 5062 757 5096
rect 757 5062 766 5096
rect 714 5053 766 5062
rect 786 5096 838 5105
rect 786 5062 795 5096
rect 795 5062 829 5096
rect 829 5062 838 5096
rect 786 5053 838 5062
rect 972 5096 1024 5105
rect 972 5062 981 5096
rect 981 5062 1015 5096
rect 1015 5062 1024 5096
rect 972 5053 1024 5062
rect 1044 5096 1096 5105
rect 1044 5062 1053 5096
rect 1053 5062 1087 5096
rect 1087 5062 1096 5096
rect 1044 5053 1096 5062
rect 198 4786 250 4795
rect 198 4752 207 4786
rect 207 4752 241 4786
rect 241 4752 250 4786
rect 198 4743 250 4752
rect 270 4786 322 4795
rect 270 4752 279 4786
rect 279 4752 313 4786
rect 313 4752 322 4786
rect 270 4743 322 4752
rect 456 4786 508 4795
rect 456 4752 465 4786
rect 465 4752 499 4786
rect 499 4752 508 4786
rect 456 4743 508 4752
rect 528 4786 580 4795
rect 528 4752 537 4786
rect 537 4752 571 4786
rect 571 4752 580 4786
rect 528 4743 580 4752
rect 198 4678 250 4687
rect 198 4644 207 4678
rect 207 4644 241 4678
rect 241 4644 250 4678
rect 198 4635 250 4644
rect 270 4678 322 4687
rect 270 4644 279 4678
rect 279 4644 313 4678
rect 313 4644 322 4678
rect 270 4635 322 4644
rect 456 4678 508 4687
rect 456 4644 465 4678
rect 465 4644 499 4678
rect 499 4644 508 4678
rect 456 4635 508 4644
rect 528 4678 580 4687
rect 528 4644 537 4678
rect 537 4644 571 4678
rect 571 4644 580 4678
rect 528 4635 580 4644
rect -318 4368 -266 4377
rect -318 4334 -309 4368
rect -309 4334 -275 4368
rect -275 4334 -266 4368
rect -318 4325 -266 4334
rect -246 4368 -194 4377
rect -246 4334 -237 4368
rect -237 4334 -203 4368
rect -203 4334 -194 4368
rect -246 4325 -194 4334
rect -60 4368 -8 4377
rect -60 4334 -51 4368
rect -51 4334 -17 4368
rect -17 4334 -8 4368
rect -60 4325 -8 4334
rect 12 4368 64 4377
rect 12 4334 21 4368
rect 21 4334 55 4368
rect 55 4334 64 4368
rect 12 4325 64 4334
rect -318 4260 -266 4269
rect -318 4226 -309 4260
rect -309 4226 -275 4260
rect -275 4226 -266 4260
rect -318 4217 -266 4226
rect -246 4260 -194 4269
rect -246 4226 -237 4260
rect -237 4226 -203 4260
rect -203 4226 -194 4260
rect -246 4217 -194 4226
rect -60 4260 -8 4269
rect -60 4226 -51 4260
rect -51 4226 -17 4260
rect -17 4226 -8 4260
rect -60 4217 -8 4226
rect 12 4260 64 4269
rect 12 4226 21 4260
rect 21 4226 55 4260
rect 55 4226 64 4260
rect 12 4217 64 4226
rect -153 4141 -101 4150
rect -153 4107 -144 4141
rect -144 4107 -110 4141
rect -110 4107 -101 4141
rect -153 4098 -101 4107
rect -153 4069 -101 4078
rect -153 4035 -144 4069
rect -144 4035 -110 4069
rect -110 4035 -101 4069
rect -153 4026 -101 4035
rect 363 4559 415 4568
rect 363 4525 372 4559
rect 372 4525 406 4559
rect 406 4525 415 4559
rect 363 4516 415 4525
rect 363 4487 415 4496
rect 363 4453 372 4487
rect 372 4453 406 4487
rect 406 4453 415 4487
rect 363 4444 415 4453
rect 879 4977 931 4986
rect 879 4943 888 4977
rect 888 4943 922 4977
rect 922 4943 931 4977
rect 879 4934 931 4943
rect 879 4905 931 4914
rect 879 4871 888 4905
rect 888 4871 922 4905
rect 922 4871 931 4905
rect 879 4862 931 4871
rect 3964 7383 4016 7392
rect 3964 7349 3973 7383
rect 3973 7349 4007 7383
rect 4007 7349 4016 7383
rect 3964 7340 4016 7349
rect 4036 7383 4088 7392
rect 4036 7349 4045 7383
rect 4045 7349 4079 7383
rect 4079 7349 4088 7383
rect 4036 7340 4088 7349
rect 4222 7383 4274 7392
rect 4222 7349 4231 7383
rect 4231 7349 4265 7383
rect 4265 7349 4274 7383
rect 4222 7340 4274 7349
rect 4294 7383 4346 7392
rect 4294 7349 4303 7383
rect 4303 7349 4337 7383
rect 4337 7349 4346 7383
rect 4294 7340 4346 7349
rect 4480 7383 4532 7392
rect 4480 7349 4489 7383
rect 4489 7349 4523 7383
rect 4523 7349 4532 7383
rect 4480 7340 4532 7349
rect 4552 7383 4604 7392
rect 4552 7349 4561 7383
rect 4561 7349 4595 7383
rect 4595 7349 4604 7383
rect 4552 7340 4604 7349
rect 4738 7383 4790 7392
rect 4738 7349 4747 7383
rect 4747 7349 4781 7383
rect 4781 7349 4790 7383
rect 4738 7340 4790 7349
rect 4810 7383 4862 7392
rect 4810 7349 4819 7383
rect 4819 7349 4853 7383
rect 4853 7349 4862 7383
rect 4810 7340 4862 7349
rect 4996 7383 5048 7392
rect 4996 7349 5005 7383
rect 5005 7349 5039 7383
rect 5039 7349 5048 7383
rect 4996 7340 5048 7349
rect 5068 7383 5120 7392
rect 5068 7349 5077 7383
rect 5077 7349 5111 7383
rect 5111 7349 5120 7383
rect 5068 7340 5120 7349
rect 5254 7383 5306 7392
rect 5254 7349 5263 7383
rect 5263 7349 5297 7383
rect 5297 7349 5306 7383
rect 5254 7340 5306 7349
rect 5326 7383 5378 7392
rect 5326 7349 5335 7383
rect 5335 7349 5369 7383
rect 5369 7349 5378 7383
rect 5326 7340 5378 7349
rect 5512 7383 5564 7392
rect 5512 7349 5521 7383
rect 5521 7349 5555 7383
rect 5555 7349 5564 7383
rect 5512 7340 5564 7349
rect 5584 7383 5636 7392
rect 5584 7349 5593 7383
rect 5593 7349 5627 7383
rect 5627 7349 5636 7383
rect 5584 7340 5636 7349
rect 5770 7383 5822 7392
rect 5770 7349 5779 7383
rect 5779 7349 5813 7383
rect 5813 7349 5822 7383
rect 5770 7340 5822 7349
rect 5842 7383 5894 7392
rect 5842 7349 5851 7383
rect 5851 7349 5885 7383
rect 5885 7349 5894 7383
rect 5842 7340 5894 7349
rect 4129 7264 4181 7273
rect 4129 7230 4138 7264
rect 4138 7230 4172 7264
rect 4172 7230 4181 7264
rect 4129 7221 4181 7230
rect 4129 7192 4181 7201
rect 4129 7158 4138 7192
rect 4138 7158 4172 7192
rect 4172 7158 4181 7192
rect 4129 7149 4181 7158
rect 3964 6965 4016 6974
rect 3964 6931 3973 6965
rect 3973 6931 4007 6965
rect 4007 6931 4016 6965
rect 3964 6922 4016 6931
rect 4036 6965 4088 6974
rect 4036 6931 4045 6965
rect 4045 6931 4079 6965
rect 4079 6931 4088 6965
rect 4036 6922 4088 6931
rect 4222 6965 4274 6974
rect 4222 6931 4231 6965
rect 4231 6931 4265 6965
rect 4265 6931 4274 6965
rect 4222 6922 4274 6931
rect 4294 6965 4346 6974
rect 4294 6931 4303 6965
rect 4303 6931 4337 6965
rect 4337 6931 4346 6965
rect 4294 6922 4346 6931
rect 4129 6846 4181 6855
rect 4129 6812 4138 6846
rect 4138 6812 4172 6846
rect 4172 6812 4181 6846
rect 4129 6803 4181 6812
rect 4129 6774 4181 6783
rect 4129 6740 4138 6774
rect 4138 6740 4172 6774
rect 4172 6740 4181 6774
rect 4129 6731 4181 6740
rect 4645 7264 4697 7273
rect 4645 7230 4654 7264
rect 4654 7230 4688 7264
rect 4688 7230 4697 7264
rect 4645 7221 4697 7230
rect 4645 7192 4697 7201
rect 4645 7158 4654 7192
rect 4654 7158 4688 7192
rect 4688 7158 4697 7192
rect 4645 7149 4697 7158
rect 4129 6428 4181 6437
rect 4129 6394 4138 6428
rect 4138 6394 4172 6428
rect 4172 6394 4181 6428
rect 4129 6385 4181 6394
rect 4129 6356 4181 6365
rect 4129 6322 4138 6356
rect 4138 6322 4172 6356
rect 4172 6322 4181 6356
rect 4129 6313 4181 6322
rect 4645 6846 4697 6855
rect 4645 6812 4654 6846
rect 4654 6812 4688 6846
rect 4688 6812 4697 6846
rect 4645 6803 4697 6812
rect 4645 6774 4697 6783
rect 4645 6740 4654 6774
rect 4654 6740 4688 6774
rect 4688 6740 4697 6774
rect 4645 6731 4697 6740
rect 5161 7264 5213 7273
rect 5161 7230 5170 7264
rect 5170 7230 5204 7264
rect 5204 7230 5213 7264
rect 5161 7221 5213 7230
rect 5161 7192 5213 7201
rect 5161 7158 5170 7192
rect 5170 7158 5204 7192
rect 5204 7158 5213 7192
rect 5161 7149 5213 7158
rect 4996 6965 5048 6974
rect 4996 6931 5005 6965
rect 5005 6931 5039 6965
rect 5039 6931 5048 6965
rect 4996 6922 5048 6931
rect 5068 6965 5120 6974
rect 5068 6931 5077 6965
rect 5077 6931 5111 6965
rect 5111 6931 5120 6965
rect 5068 6922 5120 6931
rect 5254 6965 5306 6974
rect 5254 6931 5263 6965
rect 5263 6931 5297 6965
rect 5297 6931 5306 6965
rect 5254 6922 5306 6931
rect 5326 6965 5378 6974
rect 5326 6931 5335 6965
rect 5335 6931 5369 6965
rect 5369 6931 5378 6965
rect 5326 6922 5378 6931
rect 4480 6655 4532 6664
rect 4480 6621 4489 6655
rect 4489 6621 4523 6655
rect 4523 6621 4532 6655
rect 4480 6612 4532 6621
rect 4552 6655 4604 6664
rect 4552 6621 4561 6655
rect 4561 6621 4595 6655
rect 4595 6621 4604 6655
rect 4552 6612 4604 6621
rect 4738 6655 4790 6664
rect 4738 6621 4747 6655
rect 4747 6621 4781 6655
rect 4781 6621 4790 6655
rect 4738 6612 4790 6621
rect 4810 6655 4862 6664
rect 4810 6621 4819 6655
rect 4819 6621 4853 6655
rect 4853 6621 4862 6655
rect 4810 6612 4862 6621
rect 4480 6547 4532 6556
rect 4480 6513 4489 6547
rect 4489 6513 4523 6547
rect 4523 6513 4532 6547
rect 4480 6504 4532 6513
rect 4552 6547 4604 6556
rect 4552 6513 4561 6547
rect 4561 6513 4595 6547
rect 4595 6513 4604 6547
rect 4552 6504 4604 6513
rect 4738 6547 4790 6556
rect 4738 6513 4747 6547
rect 4747 6513 4781 6547
rect 4781 6513 4790 6547
rect 4738 6504 4790 6513
rect 4810 6547 4862 6556
rect 4810 6513 4819 6547
rect 4819 6513 4853 6547
rect 4853 6513 4862 6547
rect 4810 6504 4862 6513
rect 3964 6237 4016 6246
rect 3964 6203 3973 6237
rect 3973 6203 4007 6237
rect 4007 6203 4016 6237
rect 3964 6194 4016 6203
rect 4036 6237 4088 6246
rect 4036 6203 4045 6237
rect 4045 6203 4079 6237
rect 4079 6203 4088 6237
rect 4036 6194 4088 6203
rect 4222 6237 4274 6246
rect 4222 6203 4231 6237
rect 4231 6203 4265 6237
rect 4265 6203 4274 6237
rect 4222 6194 4274 6203
rect 4294 6237 4346 6246
rect 4294 6203 4303 6237
rect 4303 6203 4337 6237
rect 4337 6203 4346 6237
rect 4294 6194 4346 6203
rect 3964 6129 4016 6138
rect 3964 6095 3973 6129
rect 3973 6095 4007 6129
rect 4007 6095 4016 6129
rect 3964 6086 4016 6095
rect 4036 6129 4088 6138
rect 4036 6095 4045 6129
rect 4045 6095 4079 6129
rect 4079 6095 4088 6129
rect 4036 6086 4088 6095
rect 4222 6129 4274 6138
rect 4222 6095 4231 6129
rect 4231 6095 4265 6129
rect 4265 6095 4274 6129
rect 4222 6086 4274 6095
rect 4294 6129 4346 6138
rect 4294 6095 4303 6129
rect 4303 6095 4337 6129
rect 4337 6095 4346 6129
rect 4294 6086 4346 6095
rect 4129 6010 4181 6019
rect 4129 5976 4138 6010
rect 4138 5976 4172 6010
rect 4172 5976 4181 6010
rect 4129 5967 4181 5976
rect 4129 5938 4181 5947
rect 4129 5904 4138 5938
rect 4138 5904 4172 5938
rect 4172 5904 4181 5938
rect 4129 5895 4181 5904
rect 4645 6428 4697 6437
rect 4645 6394 4654 6428
rect 4654 6394 4688 6428
rect 4688 6394 4697 6428
rect 4645 6385 4697 6394
rect 4645 6356 4697 6365
rect 4645 6322 4654 6356
rect 4654 6322 4688 6356
rect 4688 6322 4697 6356
rect 4645 6313 4697 6322
rect 5161 6846 5213 6855
rect 5161 6812 5170 6846
rect 5170 6812 5204 6846
rect 5204 6812 5213 6846
rect 5161 6803 5213 6812
rect 5161 6774 5213 6783
rect 5161 6740 5170 6774
rect 5170 6740 5204 6774
rect 5204 6740 5213 6774
rect 5161 6731 5213 6740
rect 5677 7264 5729 7273
rect 5677 7230 5686 7264
rect 5686 7230 5720 7264
rect 5720 7230 5729 7264
rect 5677 7221 5729 7230
rect 5677 7192 5729 7201
rect 5677 7158 5686 7192
rect 5686 7158 5720 7192
rect 5720 7158 5729 7192
rect 5677 7149 5729 7158
rect 4129 5592 4181 5601
rect 4129 5558 4138 5592
rect 4138 5558 4172 5592
rect 4172 5558 4181 5592
rect 4129 5549 4181 5558
rect 4129 5520 4181 5529
rect 4129 5486 4138 5520
rect 4138 5486 4172 5520
rect 4172 5486 4181 5520
rect 4129 5477 4181 5486
rect 4645 6010 4697 6019
rect 4645 5976 4654 6010
rect 4654 5976 4688 6010
rect 4688 5976 4697 6010
rect 4645 5967 4697 5976
rect 4645 5938 4697 5947
rect 4645 5904 4654 5938
rect 4654 5904 4688 5938
rect 4688 5904 4697 5938
rect 4645 5895 4697 5904
rect 5161 6428 5213 6437
rect 5161 6394 5170 6428
rect 5170 6394 5204 6428
rect 5204 6394 5213 6428
rect 5161 6385 5213 6394
rect 5161 6356 5213 6365
rect 5161 6322 5170 6356
rect 5170 6322 5204 6356
rect 5204 6322 5213 6356
rect 5161 6313 5213 6322
rect 5677 6846 5729 6855
rect 5677 6812 5686 6846
rect 5686 6812 5720 6846
rect 5720 6812 5729 6846
rect 5677 6803 5729 6812
rect 5677 6774 5729 6783
rect 5677 6740 5686 6774
rect 5686 6740 5720 6774
rect 5720 6740 5729 6774
rect 5677 6731 5729 6740
rect 5512 6655 5564 6664
rect 5512 6621 5521 6655
rect 5521 6621 5555 6655
rect 5555 6621 5564 6655
rect 5512 6612 5564 6621
rect 5584 6655 5636 6664
rect 5584 6621 5593 6655
rect 5593 6621 5627 6655
rect 5627 6621 5636 6655
rect 5584 6612 5636 6621
rect 5770 6655 5822 6664
rect 5770 6621 5779 6655
rect 5779 6621 5813 6655
rect 5813 6621 5822 6655
rect 5770 6612 5822 6621
rect 5842 6655 5894 6664
rect 5842 6621 5851 6655
rect 5851 6621 5885 6655
rect 5885 6621 5894 6655
rect 5842 6612 5894 6621
rect 5512 6547 5564 6556
rect 5512 6513 5521 6547
rect 5521 6513 5555 6547
rect 5555 6513 5564 6547
rect 5512 6504 5564 6513
rect 5584 6547 5636 6556
rect 5584 6513 5593 6547
rect 5593 6513 5627 6547
rect 5627 6513 5636 6547
rect 5584 6504 5636 6513
rect 5770 6547 5822 6556
rect 5770 6513 5779 6547
rect 5779 6513 5813 6547
rect 5813 6513 5822 6547
rect 5770 6504 5822 6513
rect 5842 6547 5894 6556
rect 5842 6513 5851 6547
rect 5851 6513 5885 6547
rect 5885 6513 5894 6547
rect 5842 6504 5894 6513
rect 4996 6237 5048 6246
rect 4996 6203 5005 6237
rect 5005 6203 5039 6237
rect 5039 6203 5048 6237
rect 4996 6194 5048 6203
rect 5068 6237 5120 6246
rect 5068 6203 5077 6237
rect 5077 6203 5111 6237
rect 5111 6203 5120 6237
rect 5068 6194 5120 6203
rect 5254 6237 5306 6246
rect 5254 6203 5263 6237
rect 5263 6203 5297 6237
rect 5297 6203 5306 6237
rect 5254 6194 5306 6203
rect 5326 6237 5378 6246
rect 5326 6203 5335 6237
rect 5335 6203 5369 6237
rect 5369 6203 5378 6237
rect 5326 6194 5378 6203
rect 4996 6129 5048 6138
rect 4996 6095 5005 6129
rect 5005 6095 5039 6129
rect 5039 6095 5048 6129
rect 4996 6086 5048 6095
rect 5068 6129 5120 6138
rect 5068 6095 5077 6129
rect 5077 6095 5111 6129
rect 5111 6095 5120 6129
rect 5068 6086 5120 6095
rect 5254 6129 5306 6138
rect 5254 6095 5263 6129
rect 5263 6095 5297 6129
rect 5297 6095 5306 6129
rect 5254 6086 5306 6095
rect 5326 6129 5378 6138
rect 5326 6095 5335 6129
rect 5335 6095 5369 6129
rect 5369 6095 5378 6129
rect 5326 6086 5378 6095
rect 4480 5819 4532 5828
rect 4480 5785 4489 5819
rect 4489 5785 4523 5819
rect 4523 5785 4532 5819
rect 4480 5776 4532 5785
rect 4552 5819 4604 5828
rect 4552 5785 4561 5819
rect 4561 5785 4595 5819
rect 4595 5785 4604 5819
rect 4552 5776 4604 5785
rect 4738 5819 4790 5828
rect 4738 5785 4747 5819
rect 4747 5785 4781 5819
rect 4781 5785 4790 5819
rect 4738 5776 4790 5785
rect 4810 5819 4862 5828
rect 4810 5785 4819 5819
rect 4819 5785 4853 5819
rect 4853 5785 4862 5819
rect 4810 5776 4862 5785
rect 4480 5711 4532 5720
rect 4480 5677 4489 5711
rect 4489 5677 4523 5711
rect 4523 5677 4532 5711
rect 4480 5668 4532 5677
rect 4552 5711 4604 5720
rect 4552 5677 4561 5711
rect 4561 5677 4595 5711
rect 4595 5677 4604 5711
rect 4552 5668 4604 5677
rect 4738 5711 4790 5720
rect 4738 5677 4747 5711
rect 4747 5677 4781 5711
rect 4781 5677 4790 5711
rect 4738 5668 4790 5677
rect 4810 5711 4862 5720
rect 4810 5677 4819 5711
rect 4819 5677 4853 5711
rect 4853 5677 4862 5711
rect 4810 5668 4862 5677
rect 3964 5401 4016 5410
rect 3964 5367 3973 5401
rect 3973 5367 4007 5401
rect 4007 5367 4016 5401
rect 3964 5358 4016 5367
rect 4036 5401 4088 5410
rect 4036 5367 4045 5401
rect 4045 5367 4079 5401
rect 4079 5367 4088 5401
rect 4036 5358 4088 5367
rect 4222 5401 4274 5410
rect 4222 5367 4231 5401
rect 4231 5367 4265 5401
rect 4265 5367 4274 5401
rect 4222 5358 4274 5367
rect 4294 5401 4346 5410
rect 4294 5367 4303 5401
rect 4303 5367 4337 5401
rect 4337 5367 4346 5401
rect 4294 5358 4346 5367
rect 3964 5293 4016 5302
rect 3964 5259 3973 5293
rect 3973 5259 4007 5293
rect 4007 5259 4016 5293
rect 3964 5250 4016 5259
rect 4036 5293 4088 5302
rect 4036 5259 4045 5293
rect 4045 5259 4079 5293
rect 4079 5259 4088 5293
rect 4036 5250 4088 5259
rect 4222 5293 4274 5302
rect 4222 5259 4231 5293
rect 4231 5259 4265 5293
rect 4265 5259 4274 5293
rect 4222 5250 4274 5259
rect 4294 5293 4346 5302
rect 4294 5259 4303 5293
rect 4303 5259 4337 5293
rect 4337 5259 4346 5293
rect 4294 5250 4346 5259
rect 4129 5174 4181 5183
rect 4129 5140 4138 5174
rect 4138 5140 4172 5174
rect 4172 5140 4181 5174
rect 4129 5131 4181 5140
rect 4129 5102 4181 5111
rect 4129 5068 4138 5102
rect 4138 5068 4172 5102
rect 4172 5068 4181 5102
rect 4129 5059 4181 5068
rect 4645 5592 4697 5601
rect 4645 5558 4654 5592
rect 4654 5558 4688 5592
rect 4688 5558 4697 5592
rect 4645 5549 4697 5558
rect 4645 5520 4697 5529
rect 4645 5486 4654 5520
rect 4654 5486 4688 5520
rect 4688 5486 4697 5520
rect 4645 5477 4697 5486
rect 5161 6010 5213 6019
rect 5161 5976 5170 6010
rect 5170 5976 5204 6010
rect 5204 5976 5213 6010
rect 5161 5967 5213 5976
rect 5161 5938 5213 5947
rect 5161 5904 5170 5938
rect 5170 5904 5204 5938
rect 5204 5904 5213 5938
rect 5161 5895 5213 5904
rect 5677 6428 5729 6437
rect 5677 6394 5686 6428
rect 5686 6394 5720 6428
rect 5720 6394 5729 6428
rect 5677 6385 5729 6394
rect 5677 6356 5729 6365
rect 5677 6322 5686 6356
rect 5686 6322 5720 6356
rect 5720 6322 5729 6356
rect 5677 6313 5729 6322
rect 4129 4756 4181 4765
rect 4129 4722 4138 4756
rect 4138 4722 4172 4756
rect 4172 4722 4181 4756
rect 4129 4713 4181 4722
rect 4129 4684 4181 4693
rect 4129 4650 4138 4684
rect 4138 4650 4172 4684
rect 4172 4650 4181 4684
rect 4129 4641 4181 4650
rect 4645 5174 4697 5183
rect 4645 5140 4654 5174
rect 4654 5140 4688 5174
rect 4688 5140 4697 5174
rect 4645 5131 4697 5140
rect 4645 5102 4697 5111
rect 4645 5068 4654 5102
rect 4654 5068 4688 5102
rect 4688 5068 4697 5102
rect 4645 5059 4697 5068
rect 5161 5592 5213 5601
rect 5161 5558 5170 5592
rect 5170 5558 5204 5592
rect 5204 5558 5213 5592
rect 5161 5549 5213 5558
rect 5161 5520 5213 5529
rect 5161 5486 5170 5520
rect 5170 5486 5204 5520
rect 5204 5486 5213 5520
rect 5161 5477 5213 5486
rect 5677 6010 5729 6019
rect 5677 5976 5686 6010
rect 5686 5976 5720 6010
rect 5720 5976 5729 6010
rect 5677 5967 5729 5976
rect 5677 5938 5729 5947
rect 5677 5904 5686 5938
rect 5686 5904 5720 5938
rect 5720 5904 5729 5938
rect 5677 5895 5729 5904
rect 5512 5819 5564 5828
rect 5512 5785 5521 5819
rect 5521 5785 5555 5819
rect 5555 5785 5564 5819
rect 5512 5776 5564 5785
rect 5584 5819 5636 5828
rect 5584 5785 5593 5819
rect 5593 5785 5627 5819
rect 5627 5785 5636 5819
rect 5584 5776 5636 5785
rect 5770 5819 5822 5828
rect 5770 5785 5779 5819
rect 5779 5785 5813 5819
rect 5813 5785 5822 5819
rect 5770 5776 5822 5785
rect 5842 5819 5894 5828
rect 5842 5785 5851 5819
rect 5851 5785 5885 5819
rect 5885 5785 5894 5819
rect 5842 5776 5894 5785
rect 5512 5711 5564 5720
rect 5512 5677 5521 5711
rect 5521 5677 5555 5711
rect 5555 5677 5564 5711
rect 5512 5668 5564 5677
rect 5584 5711 5636 5720
rect 5584 5677 5593 5711
rect 5593 5677 5627 5711
rect 5627 5677 5636 5711
rect 5584 5668 5636 5677
rect 5770 5711 5822 5720
rect 5770 5677 5779 5711
rect 5779 5677 5813 5711
rect 5813 5677 5822 5711
rect 5770 5668 5822 5677
rect 5842 5711 5894 5720
rect 5842 5677 5851 5711
rect 5851 5677 5885 5711
rect 5885 5677 5894 5711
rect 5842 5668 5894 5677
rect 4996 5401 5048 5410
rect 4996 5367 5005 5401
rect 5005 5367 5039 5401
rect 5039 5367 5048 5401
rect 4996 5358 5048 5367
rect 5068 5401 5120 5410
rect 5068 5367 5077 5401
rect 5077 5367 5111 5401
rect 5111 5367 5120 5401
rect 5068 5358 5120 5367
rect 5254 5401 5306 5410
rect 5254 5367 5263 5401
rect 5263 5367 5297 5401
rect 5297 5367 5306 5401
rect 5254 5358 5306 5367
rect 5326 5401 5378 5410
rect 5326 5367 5335 5401
rect 5335 5367 5369 5401
rect 5369 5367 5378 5401
rect 5326 5358 5378 5367
rect 4996 5293 5048 5302
rect 4996 5259 5005 5293
rect 5005 5259 5039 5293
rect 5039 5259 5048 5293
rect 4996 5250 5048 5259
rect 5068 5293 5120 5302
rect 5068 5259 5077 5293
rect 5077 5259 5111 5293
rect 5111 5259 5120 5293
rect 5068 5250 5120 5259
rect 5254 5293 5306 5302
rect 5254 5259 5263 5293
rect 5263 5259 5297 5293
rect 5297 5259 5306 5293
rect 5254 5250 5306 5259
rect 5326 5293 5378 5302
rect 5326 5259 5335 5293
rect 5335 5259 5369 5293
rect 5369 5259 5378 5293
rect 5326 5250 5378 5259
rect 4480 4983 4532 4992
rect 4480 4949 4489 4983
rect 4489 4949 4523 4983
rect 4523 4949 4532 4983
rect 4480 4940 4532 4949
rect 4552 4983 4604 4992
rect 4552 4949 4561 4983
rect 4561 4949 4595 4983
rect 4595 4949 4604 4983
rect 4552 4940 4604 4949
rect 4738 4983 4790 4992
rect 4738 4949 4747 4983
rect 4747 4949 4781 4983
rect 4781 4949 4790 4983
rect 4738 4940 4790 4949
rect 4810 4983 4862 4992
rect 4810 4949 4819 4983
rect 4819 4949 4853 4983
rect 4853 4949 4862 4983
rect 4810 4940 4862 4949
rect 4480 4875 4532 4884
rect 4480 4841 4489 4875
rect 4489 4841 4523 4875
rect 4523 4841 4532 4875
rect 4480 4832 4532 4841
rect 4552 4875 4604 4884
rect 4552 4841 4561 4875
rect 4561 4841 4595 4875
rect 4595 4841 4604 4875
rect 4552 4832 4604 4841
rect 4738 4875 4790 4884
rect 4738 4841 4747 4875
rect 4747 4841 4781 4875
rect 4781 4841 4790 4875
rect 4738 4832 4790 4841
rect 4810 4875 4862 4884
rect 4810 4841 4819 4875
rect 4819 4841 4853 4875
rect 4853 4841 4862 4875
rect 4810 4832 4862 4841
rect 3964 4565 4016 4574
rect 3964 4531 3973 4565
rect 3973 4531 4007 4565
rect 4007 4531 4016 4565
rect 3964 4522 4016 4531
rect 4036 4565 4088 4574
rect 4036 4531 4045 4565
rect 4045 4531 4079 4565
rect 4079 4531 4088 4565
rect 4036 4522 4088 4531
rect 4222 4565 4274 4574
rect 4222 4531 4231 4565
rect 4231 4531 4265 4565
rect 4265 4531 4274 4565
rect 4222 4522 4274 4531
rect 4294 4565 4346 4574
rect 4294 4531 4303 4565
rect 4303 4531 4337 4565
rect 4337 4531 4346 4565
rect 4294 4522 4346 4531
rect 3964 4457 4016 4466
rect 3964 4423 3973 4457
rect 3973 4423 4007 4457
rect 4007 4423 4016 4457
rect 3964 4414 4016 4423
rect 4036 4457 4088 4466
rect 4036 4423 4045 4457
rect 4045 4423 4079 4457
rect 4079 4423 4088 4457
rect 4036 4414 4088 4423
rect 4222 4457 4274 4466
rect 4222 4423 4231 4457
rect 4231 4423 4265 4457
rect 4265 4423 4274 4457
rect 4222 4414 4274 4423
rect 4294 4457 4346 4466
rect 4294 4423 4303 4457
rect 4303 4423 4337 4457
rect 4337 4423 4346 4457
rect 4294 4414 4346 4423
rect 1395 4035 1404 4050
rect 1404 4035 1438 4050
rect 1438 4035 1447 4050
rect 1395 3998 1447 4035
rect 1509 4041 1561 4050
rect 1509 4007 1518 4041
rect 1518 4007 1552 4041
rect 1552 4007 1561 4041
rect 1509 3998 1561 4007
rect 4129 4338 4181 4347
rect 4129 4304 4138 4338
rect 4138 4304 4172 4338
rect 4172 4304 4181 4338
rect 4129 4295 4181 4304
rect 4129 4266 4181 4275
rect 4129 4232 4138 4266
rect 4138 4232 4172 4266
rect 4172 4232 4181 4266
rect 4129 4223 4181 4232
rect 4645 4756 4697 4765
rect 4645 4722 4654 4756
rect 4654 4722 4688 4756
rect 4688 4722 4697 4756
rect 4645 4713 4697 4722
rect 4645 4684 4697 4693
rect 4645 4650 4654 4684
rect 4654 4650 4688 4684
rect 4688 4650 4697 4684
rect 4645 4641 4697 4650
rect 5161 5174 5213 5183
rect 5161 5140 5170 5174
rect 5170 5140 5204 5174
rect 5204 5140 5213 5174
rect 5161 5131 5213 5140
rect 5161 5102 5213 5111
rect 5161 5068 5170 5102
rect 5170 5068 5204 5102
rect 5204 5068 5213 5102
rect 5161 5059 5213 5068
rect 5677 5592 5729 5601
rect 5677 5558 5686 5592
rect 5686 5558 5720 5592
rect 5720 5558 5729 5592
rect 5677 5549 5729 5558
rect 5677 5520 5729 5529
rect 5677 5486 5686 5520
rect 5686 5486 5720 5520
rect 5720 5486 5729 5520
rect 5677 5477 5729 5486
rect 4480 4457 4532 4466
rect 4480 4423 4489 4457
rect 4489 4423 4523 4457
rect 4523 4423 4532 4457
rect 4480 4414 4532 4423
rect 4552 4457 4604 4466
rect 4552 4423 4561 4457
rect 4561 4423 4595 4457
rect 4595 4423 4604 4457
rect 4552 4414 4604 4423
rect 4738 4457 4790 4466
rect 4738 4423 4747 4457
rect 4747 4423 4781 4457
rect 4781 4423 4790 4457
rect 4738 4414 4790 4423
rect 4810 4457 4862 4466
rect 4810 4423 4819 4457
rect 4819 4423 4853 4457
rect 4853 4423 4862 4457
rect 4810 4414 4862 4423
rect 4645 4338 4697 4347
rect 4645 4304 4654 4338
rect 4654 4304 4688 4338
rect 4688 4304 4697 4338
rect 4645 4295 4697 4304
rect 4645 4266 4697 4275
rect 4645 4232 4654 4266
rect 4654 4232 4688 4266
rect 4688 4232 4697 4266
rect 4645 4223 4697 4232
rect 5161 4756 5213 4765
rect 5161 4722 5170 4756
rect 5170 4722 5204 4756
rect 5204 4722 5213 4756
rect 5161 4713 5213 4722
rect 5161 4684 5213 4693
rect 5161 4650 5170 4684
rect 5170 4650 5204 4684
rect 5204 4650 5213 4684
rect 5161 4641 5213 4650
rect 5677 5174 5729 5183
rect 5677 5140 5686 5174
rect 5686 5140 5720 5174
rect 5720 5140 5729 5174
rect 5677 5131 5729 5140
rect 5677 5102 5729 5111
rect 5677 5068 5686 5102
rect 5686 5068 5720 5102
rect 5720 5068 5729 5102
rect 5677 5059 5729 5068
rect 5512 4983 5564 4992
rect 5512 4949 5521 4983
rect 5521 4949 5555 4983
rect 5555 4949 5564 4983
rect 5512 4940 5564 4949
rect 5584 4983 5636 4992
rect 5584 4949 5593 4983
rect 5593 4949 5627 4983
rect 5627 4949 5636 4983
rect 5584 4940 5636 4949
rect 5770 4983 5822 4992
rect 5770 4949 5779 4983
rect 5779 4949 5813 4983
rect 5813 4949 5822 4983
rect 5770 4940 5822 4949
rect 5842 4983 5894 4992
rect 5842 4949 5851 4983
rect 5851 4949 5885 4983
rect 5885 4949 5894 4983
rect 5842 4940 5894 4949
rect 5512 4875 5564 4884
rect 5512 4841 5521 4875
rect 5521 4841 5555 4875
rect 5555 4841 5564 4875
rect 5512 4832 5564 4841
rect 5584 4875 5636 4884
rect 5584 4841 5593 4875
rect 5593 4841 5627 4875
rect 5627 4841 5636 4875
rect 5584 4832 5636 4841
rect 5770 4875 5822 4884
rect 5770 4841 5779 4875
rect 5779 4841 5813 4875
rect 5813 4841 5822 4875
rect 5770 4832 5822 4841
rect 5842 4875 5894 4884
rect 5842 4841 5851 4875
rect 5851 4841 5885 4875
rect 5885 4841 5894 4875
rect 5842 4832 5894 4841
rect 4996 4565 5048 4574
rect 4996 4531 5005 4565
rect 5005 4531 5039 4565
rect 5039 4531 5048 4565
rect 4996 4522 5048 4531
rect 5068 4565 5120 4574
rect 5068 4531 5077 4565
rect 5077 4531 5111 4565
rect 5111 4531 5120 4565
rect 5068 4522 5120 4531
rect 5254 4565 5306 4574
rect 5254 4531 5263 4565
rect 5263 4531 5297 4565
rect 5297 4531 5306 4565
rect 5254 4522 5306 4531
rect 5326 4565 5378 4574
rect 5326 4531 5335 4565
rect 5335 4531 5369 4565
rect 5369 4531 5378 4565
rect 5326 4522 5378 4531
rect 4996 4457 5048 4466
rect 4996 4423 5005 4457
rect 5005 4423 5039 4457
rect 5039 4423 5048 4457
rect 4996 4414 5048 4423
rect 5068 4457 5120 4466
rect 5068 4423 5077 4457
rect 5077 4423 5111 4457
rect 5111 4423 5120 4457
rect 5068 4414 5120 4423
rect 5254 4457 5306 4466
rect 5254 4423 5263 4457
rect 5263 4423 5297 4457
rect 5297 4423 5306 4457
rect 5254 4414 5306 4423
rect 5326 4457 5378 4466
rect 5326 4423 5335 4457
rect 5335 4423 5369 4457
rect 5369 4423 5378 4457
rect 5326 4414 5378 4423
rect 5161 4338 5213 4347
rect 5161 4304 5170 4338
rect 5170 4304 5204 4338
rect 5204 4304 5213 4338
rect 5161 4295 5213 4304
rect 5161 4266 5213 4275
rect 5161 4232 5170 4266
rect 5170 4232 5204 4266
rect 5204 4232 5213 4266
rect 5161 4223 5213 4232
rect 5677 4756 5729 4765
rect 5677 4722 5686 4756
rect 5686 4722 5720 4756
rect 5720 4722 5729 4756
rect 5677 4713 5729 4722
rect 5677 4684 5729 4693
rect 5677 4650 5686 4684
rect 5686 4650 5720 4684
rect 5720 4650 5729 4684
rect 5677 4641 5729 4650
rect 5512 4457 5564 4466
rect 5512 4423 5521 4457
rect 5521 4423 5555 4457
rect 5555 4423 5564 4457
rect 5512 4414 5564 4423
rect 5584 4457 5636 4466
rect 5584 4423 5593 4457
rect 5593 4423 5627 4457
rect 5627 4423 5636 4457
rect 5584 4414 5636 4423
rect 5770 4457 5822 4466
rect 5770 4423 5779 4457
rect 5779 4423 5813 4457
rect 5813 4423 5822 4457
rect 5770 4414 5822 4423
rect 5842 4457 5894 4466
rect 5842 4423 5851 4457
rect 5851 4423 5885 4457
rect 5885 4423 5894 4457
rect 5842 4414 5894 4423
rect 5677 4338 5729 4347
rect 5677 4304 5686 4338
rect 5686 4304 5720 4338
rect 5720 4304 5729 4338
rect 5677 4295 5729 4304
rect 5677 4266 5729 4275
rect 5677 4232 5686 4266
rect 5686 4232 5720 4266
rect 5720 4232 5729 4266
rect 5677 4223 5729 4232
rect 6307 4238 6359 4247
rect 6307 4204 6316 4238
rect 6316 4204 6350 4238
rect 6350 4204 6359 4238
rect 6307 4195 6359 4204
rect 6519 3948 6571 4000
rect -2619 3506 -2567 3558
rect -2619 3228 -2567 3280
rect 8700 6972 8752 6981
rect 8700 6938 8709 6972
rect 8709 6938 8743 6972
rect 8743 6938 8752 6972
rect 8700 6929 8752 6938
rect 8772 6972 8824 6981
rect 8772 6938 8781 6972
rect 8781 6938 8815 6972
rect 8815 6938 8824 6972
rect 8772 6929 8824 6938
rect 8607 6853 8659 6862
rect 8607 6819 8616 6853
rect 8616 6819 8650 6853
rect 8650 6819 8659 6853
rect 8607 6810 8659 6819
rect 8958 6972 9010 6981
rect 8958 6938 8967 6972
rect 8967 6938 9001 6972
rect 9001 6938 9010 6972
rect 8958 6929 9010 6938
rect 9030 6972 9082 6981
rect 9030 6938 9039 6972
rect 9039 6938 9073 6972
rect 9073 6938 9082 6972
rect 9030 6929 9082 6938
rect 9216 6972 9268 6981
rect 9216 6938 9225 6972
rect 9225 6938 9259 6972
rect 9259 6938 9268 6972
rect 9216 6929 9268 6938
rect 9288 6972 9340 6981
rect 9288 6938 9297 6972
rect 9297 6938 9331 6972
rect 9331 6938 9340 6972
rect 9288 6929 9340 6938
rect 8700 6554 8752 6563
rect 8700 6520 8709 6554
rect 8709 6520 8743 6554
rect 8743 6520 8752 6554
rect 8700 6511 8752 6520
rect 8772 6554 8824 6563
rect 8772 6520 8781 6554
rect 8781 6520 8815 6554
rect 8815 6520 8824 6554
rect 8772 6511 8824 6520
rect 9123 6853 9175 6862
rect 9123 6819 9132 6853
rect 9132 6819 9166 6853
rect 9166 6819 9175 6853
rect 9123 6810 9175 6819
rect 9474 6972 9526 6981
rect 9474 6938 9483 6972
rect 9483 6938 9517 6972
rect 9517 6938 9526 6972
rect 9474 6929 9526 6938
rect 9546 6972 9598 6981
rect 9546 6938 9555 6972
rect 9555 6938 9589 6972
rect 9589 6938 9598 6972
rect 9546 6929 9598 6938
rect 8958 6554 9010 6563
rect 8958 6520 8967 6554
rect 8967 6520 9001 6554
rect 9001 6520 9010 6554
rect 8958 6511 9010 6520
rect 9030 6554 9082 6563
rect 9030 6520 9039 6554
rect 9039 6520 9073 6554
rect 9073 6520 9082 6554
rect 9030 6511 9082 6520
rect 8700 6136 8752 6145
rect 8700 6102 8709 6136
rect 8709 6102 8743 6136
rect 8743 6102 8752 6136
rect 8700 6093 8752 6102
rect 8772 6136 8824 6145
rect 8772 6102 8781 6136
rect 8781 6102 8815 6136
rect 8815 6102 8824 6136
rect 8772 6093 8824 6102
rect 9216 6554 9268 6563
rect 9216 6520 9225 6554
rect 9225 6520 9259 6554
rect 9259 6520 9268 6554
rect 9216 6511 9268 6520
rect 9288 6554 9340 6563
rect 9288 6520 9297 6554
rect 9297 6520 9331 6554
rect 9331 6520 9340 6554
rect 9288 6511 9340 6520
rect 8958 6136 9010 6145
rect 8958 6102 8967 6136
rect 8967 6102 9001 6136
rect 9001 6102 9010 6136
rect 8958 6093 9010 6102
rect 9030 6136 9082 6145
rect 9030 6102 9039 6136
rect 9039 6102 9073 6136
rect 9073 6102 9082 6136
rect 9030 6093 9082 6102
rect 8700 5718 8752 5727
rect 8700 5684 8709 5718
rect 8709 5684 8743 5718
rect 8743 5684 8752 5718
rect 8700 5675 8752 5684
rect 8772 5718 8824 5727
rect 8772 5684 8781 5718
rect 8781 5684 8815 5718
rect 8815 5684 8824 5718
rect 8772 5675 8824 5684
rect 8607 5599 8659 5608
rect 8607 5565 8616 5599
rect 8616 5565 8650 5599
rect 8650 5565 8659 5599
rect 8607 5556 8659 5565
rect 8607 5527 8659 5536
rect 8607 5493 8616 5527
rect 8616 5493 8650 5527
rect 8650 5493 8659 5527
rect 8607 5484 8659 5493
rect 9639 6853 9691 6862
rect 9639 6819 9648 6853
rect 9648 6819 9682 6853
rect 9682 6819 9691 6853
rect 9639 6810 9691 6819
rect 9474 6554 9526 6563
rect 9474 6520 9483 6554
rect 9483 6520 9517 6554
rect 9517 6520 9526 6554
rect 9474 6511 9526 6520
rect 9546 6554 9598 6563
rect 9546 6520 9555 6554
rect 9555 6520 9589 6554
rect 9589 6520 9598 6554
rect 9546 6511 9598 6520
rect 9216 6136 9268 6145
rect 9216 6102 9225 6136
rect 9225 6102 9259 6136
rect 9259 6102 9268 6136
rect 9216 6093 9268 6102
rect 9288 6136 9340 6145
rect 9288 6102 9297 6136
rect 9297 6102 9331 6136
rect 9331 6102 9340 6136
rect 9288 6093 9340 6102
rect 9474 6136 9526 6145
rect 9474 6102 9483 6136
rect 9483 6102 9517 6136
rect 9517 6102 9526 6136
rect 9474 6093 9526 6102
rect 9546 6136 9598 6145
rect 9546 6102 9555 6136
rect 9555 6102 9589 6136
rect 9589 6102 9598 6136
rect 9546 6093 9598 6102
rect 8958 5718 9010 5727
rect 8958 5684 8967 5718
rect 8967 5684 9001 5718
rect 9001 5684 9010 5718
rect 8958 5675 9010 5684
rect 9030 5718 9082 5727
rect 9030 5684 9039 5718
rect 9039 5684 9073 5718
rect 9073 5684 9082 5718
rect 9030 5675 9082 5684
rect 9216 5718 9268 5727
rect 9216 5684 9225 5718
rect 9225 5684 9259 5718
rect 9259 5684 9268 5718
rect 9216 5675 9268 5684
rect 9288 5718 9340 5727
rect 9288 5684 9297 5718
rect 9297 5684 9331 5718
rect 9331 5684 9340 5718
rect 9288 5675 9340 5684
rect 8700 5300 8752 5309
rect 8700 5266 8709 5300
rect 8709 5266 8743 5300
rect 8743 5266 8752 5300
rect 8700 5257 8752 5266
rect 8772 5300 8824 5309
rect 8772 5266 8781 5300
rect 8781 5266 8815 5300
rect 8815 5266 8824 5300
rect 8772 5257 8824 5266
rect 9123 5599 9175 5608
rect 9123 5565 9132 5599
rect 9132 5565 9166 5599
rect 9166 5565 9175 5599
rect 9123 5556 9175 5565
rect 9123 5527 9175 5536
rect 9123 5493 9132 5527
rect 9132 5493 9166 5527
rect 9166 5493 9175 5527
rect 9123 5484 9175 5493
rect 9474 5718 9526 5727
rect 9474 5684 9483 5718
rect 9483 5684 9517 5718
rect 9517 5684 9526 5718
rect 9474 5675 9526 5684
rect 9546 5718 9598 5727
rect 9546 5684 9555 5718
rect 9555 5684 9589 5718
rect 9589 5684 9598 5718
rect 9546 5675 9598 5684
rect 8958 5300 9010 5309
rect 8958 5266 8967 5300
rect 8967 5266 9001 5300
rect 9001 5266 9010 5300
rect 8958 5257 9010 5266
rect 9030 5300 9082 5309
rect 9030 5266 9039 5300
rect 9039 5266 9073 5300
rect 9073 5266 9082 5300
rect 9030 5257 9082 5266
rect 8700 4882 8752 4891
rect 8700 4848 8709 4882
rect 8709 4848 8743 4882
rect 8743 4848 8752 4882
rect 8700 4839 8752 4848
rect 8772 4882 8824 4891
rect 8772 4848 8781 4882
rect 8781 4848 8815 4882
rect 8815 4848 8824 4882
rect 8772 4839 8824 4848
rect 9216 5300 9268 5309
rect 9216 5266 9225 5300
rect 9225 5266 9259 5300
rect 9259 5266 9268 5300
rect 9216 5257 9268 5266
rect 9288 5300 9340 5309
rect 9288 5266 9297 5300
rect 9297 5266 9331 5300
rect 9331 5266 9340 5300
rect 9288 5257 9340 5266
rect 8958 4882 9010 4891
rect 8958 4848 8967 4882
rect 8967 4848 9001 4882
rect 9001 4848 9010 4882
rect 8958 4839 9010 4848
rect 9030 4882 9082 4891
rect 9030 4848 9039 4882
rect 9039 4848 9073 4882
rect 9073 4848 9082 4882
rect 9030 4839 9082 4848
rect 8700 4464 8752 4473
rect 8700 4430 8709 4464
rect 8709 4430 8743 4464
rect 8743 4430 8752 4464
rect 8700 4421 8752 4430
rect 8772 4464 8824 4473
rect 8772 4430 8781 4464
rect 8781 4430 8815 4464
rect 8815 4430 8824 4464
rect 8772 4421 8824 4430
rect 9639 5599 9691 5608
rect 9639 5565 9648 5599
rect 9648 5565 9682 5599
rect 9682 5565 9691 5599
rect 9639 5556 9691 5565
rect 9639 5527 9691 5536
rect 9639 5493 9648 5527
rect 9648 5493 9682 5527
rect 9682 5493 9691 5527
rect 9639 5484 9691 5493
rect 9474 5300 9526 5309
rect 9474 5266 9483 5300
rect 9483 5266 9517 5300
rect 9517 5266 9526 5300
rect 9474 5257 9526 5266
rect 9546 5300 9598 5309
rect 9546 5266 9555 5300
rect 9555 5266 9589 5300
rect 9589 5266 9598 5300
rect 9546 5257 9598 5266
rect 9216 4882 9268 4891
rect 9216 4848 9225 4882
rect 9225 4848 9259 4882
rect 9259 4848 9268 4882
rect 9216 4839 9268 4848
rect 9288 4882 9340 4891
rect 9288 4848 9297 4882
rect 9297 4848 9331 4882
rect 9331 4848 9340 4882
rect 9288 4839 9340 4848
rect 8958 4464 9010 4473
rect 8958 4430 8967 4464
rect 8967 4430 9001 4464
rect 9001 4430 9010 4464
rect 8958 4421 9010 4430
rect 9030 4464 9082 4473
rect 9030 4430 9039 4464
rect 9039 4430 9073 4464
rect 9073 4430 9082 4464
rect 9030 4421 9082 4430
rect 9474 4882 9526 4891
rect 9474 4848 9483 4882
rect 9483 4848 9517 4882
rect 9517 4848 9526 4882
rect 9474 4839 9526 4848
rect 9546 4882 9598 4891
rect 9546 4848 9555 4882
rect 9555 4848 9589 4882
rect 9589 4848 9598 4882
rect 9546 4839 9598 4848
rect 9216 4464 9268 4473
rect 9216 4430 9225 4464
rect 9225 4430 9259 4464
rect 9259 4430 9268 4464
rect 9216 4421 9268 4430
rect 9288 4464 9340 4473
rect 9288 4430 9297 4464
rect 9297 4430 9331 4464
rect 9331 4430 9340 4464
rect 9288 4421 9340 4430
rect 8349 3744 8401 3796
rect 9474 4464 9526 4473
rect 9474 4430 9483 4464
rect 9483 4430 9517 4464
rect 9517 4430 9526 4464
rect 9474 4421 9526 4430
rect 9546 4464 9598 4473
rect 9546 4430 9555 4464
rect 9555 4430 9589 4464
rect 9589 4430 9598 4464
rect 9546 4421 9598 4430
rect 11107 4195 11159 4247
rect 7249 3219 7301 3271
<< metal2 >>
rect -5029 11118 5667 11164
rect -1824 10959 2818 10968
rect -1824 10903 2753 10959
rect 2809 10903 2818 10959
rect -1824 10894 2818 10903
rect -1824 10242 -1772 10894
rect 2543 10728 3683 10780
rect 3735 10728 3755 10780
rect 3807 10728 4457 10780
rect 4509 10728 4529 10780
rect 4581 10728 4615 10780
rect -227 10443 -153 10480
rect 886 10468 960 10490
rect 886 10443 895 10468
rect -227 10442 895 10443
rect -227 10390 -216 10442
rect -164 10412 895 10442
rect 951 10412 960 10468
rect -164 10391 960 10412
rect -164 10390 -153 10391
rect -227 10370 -153 10390
rect -227 10318 -216 10370
rect -164 10318 -153 10370
rect -227 10280 -153 10318
rect -1824 10190 -897 10242
rect -845 10190 -825 10242
rect -773 10190 -639 10242
rect -587 10190 -567 10242
rect -515 10190 -381 10242
rect -329 10190 -309 10242
rect -257 10190 -123 10242
rect -71 10190 -51 10242
rect 1 10190 39 10242
rect -1824 10134 -1772 10190
rect -1824 10082 -897 10134
rect -845 10082 -825 10134
rect -773 10082 -639 10134
rect -587 10082 -567 10134
rect -515 10082 -381 10134
rect -329 10082 -309 10134
rect -257 10082 -123 10134
rect -71 10082 -51 10134
rect 1 10082 39 10134
rect -1824 9370 -1772 10082
rect -743 10006 -669 10044
rect 886 10006 960 10391
rect -743 9954 -732 10006
rect -680 9954 960 10006
rect -743 9934 -669 9954
rect -743 9882 -732 9934
rect -680 9882 -669 9934
rect -743 9844 -669 9882
rect -227 9570 -153 9608
rect 886 9570 960 9954
rect -227 9518 -216 9570
rect -164 9518 960 9570
rect -227 9498 -153 9518
rect -227 9446 -216 9498
rect -164 9446 -153 9498
rect -227 9408 -153 9446
rect -1824 9318 -897 9370
rect -845 9318 -825 9370
rect -773 9318 -639 9370
rect -587 9318 -567 9370
rect -515 9318 -381 9370
rect -329 9318 -309 9370
rect -257 9318 -123 9370
rect -71 9318 -51 9370
rect 1 9318 39 9370
rect -1824 9262 -1772 9318
rect -1824 9210 -897 9262
rect -845 9210 -825 9262
rect -773 9210 -639 9262
rect -587 9210 -567 9262
rect -515 9210 -381 9262
rect -329 9210 -309 9262
rect -257 9210 -123 9262
rect -71 9210 -51 9262
rect 1 9210 39 9262
rect -1824 8837 -1772 9210
rect -743 9134 -669 9172
rect 886 9134 960 9518
rect -743 9082 -732 9134
rect -680 9082 960 9134
rect -743 9062 -669 9082
rect -743 9010 -732 9062
rect -680 9010 -669 9062
rect -743 8972 -669 9010
rect 886 8895 960 9082
rect 2543 10362 2589 10728
rect 3579 10690 3653 10699
rect 3579 10634 3588 10690
rect 3644 10634 3653 10690
rect 3579 10609 3590 10634
rect 3642 10609 3653 10634
rect 3579 10589 3653 10609
rect 3579 10537 3590 10589
rect 3642 10537 3653 10589
rect 3579 10499 3653 10537
rect 4095 10661 4169 10699
rect 4095 10609 4106 10661
rect 4158 10609 4169 10661
rect 4095 10589 4169 10609
rect 4095 10562 4106 10589
rect 4158 10562 4169 10589
rect 4095 10506 4104 10562
rect 4160 10506 4169 10562
rect 4095 10495 4169 10506
rect 4611 10690 4685 10699
rect 4611 10634 4620 10690
rect 4676 10634 4685 10690
rect 4611 10609 4622 10634
rect 4674 10609 4685 10634
rect 4611 10589 4685 10609
rect 4611 10537 4622 10589
rect 4674 10537 4685 10589
rect 4611 10499 4685 10537
rect 5621 10467 5667 11118
rect 9134 11139 9208 11148
rect 9134 11083 9143 11139
rect 9199 11083 9208 11139
rect 9134 10560 9208 11083
rect 10013 11139 10087 11148
rect 10013 11083 10022 11139
rect 10078 11083 10087 11139
rect 10013 10838 10087 11083
rect 10013 10829 10088 10838
rect 10013 10777 10024 10829
rect 10076 10777 10088 10829
rect 10013 10765 10088 10777
rect 10014 10764 10088 10765
rect 7335 10508 7351 10560
rect 7403 10508 7423 10560
rect 7475 10508 7609 10560
rect 7661 10508 7681 10560
rect 7733 10508 7867 10560
rect 7919 10508 7939 10560
rect 7991 10508 8125 10560
rect 8177 10508 8197 10560
rect 8249 10508 9208 10560
rect 3907 10415 3941 10467
rect 3993 10415 4013 10467
rect 4065 10415 4199 10467
rect 4251 10415 4271 10467
rect 4323 10415 5667 10467
rect 9134 10452 9208 10508
rect 2543 10310 3941 10362
rect 3993 10310 4013 10362
rect 4065 10310 4199 10362
rect 4251 10310 4271 10362
rect 4323 10310 4357 10362
rect 2543 9944 2589 10310
rect 3579 10243 3653 10281
rect 3579 10191 3590 10243
rect 3642 10191 3653 10243
rect 3579 10171 3653 10191
rect 3579 10142 3590 10171
rect 3642 10142 3653 10171
rect 3579 10086 3588 10142
rect 3644 10086 3653 10142
rect 3579 10077 3653 10086
rect 4095 10271 4169 10281
rect 4095 10215 4104 10271
rect 4160 10215 4169 10271
rect 4095 10191 4106 10215
rect 4158 10191 4169 10215
rect 4095 10171 4169 10191
rect 4095 10119 4106 10171
rect 4158 10119 4169 10171
rect 4095 10081 4169 10119
rect 4611 10243 4685 10281
rect 4611 10191 4622 10243
rect 4674 10191 4685 10243
rect 4611 10171 4685 10191
rect 4611 10141 4622 10171
rect 4674 10141 4685 10171
rect 4611 10085 4620 10141
rect 4676 10085 4685 10141
rect 4611 10077 4685 10085
rect 5621 10049 5667 10415
rect 7335 10400 7351 10452
rect 7403 10400 7423 10452
rect 7475 10400 7609 10452
rect 7661 10400 7681 10452
rect 7733 10400 7867 10452
rect 7919 10400 7939 10452
rect 7991 10400 8125 10452
rect 8177 10400 8197 10452
rect 8249 10400 9208 10452
rect 3391 9997 3425 10049
rect 3477 9997 3497 10049
rect 3549 9997 3683 10049
rect 3735 9997 3755 10049
rect 3807 9997 4457 10049
rect 4509 9997 4529 10049
rect 4581 9997 4715 10049
rect 4767 9997 4787 10049
rect 4839 9997 5667 10049
rect 2543 9892 3425 9944
rect 3477 9892 3497 9944
rect 3549 9892 3683 9944
rect 3735 9892 3755 9944
rect 3807 9892 4457 9944
rect 4509 9892 4529 9944
rect 4581 9892 4715 9944
rect 4767 9892 4787 9944
rect 4839 9892 4873 9944
rect 2543 9526 2589 9892
rect 3579 9854 3653 9863
rect 3579 9798 3588 9854
rect 3644 9798 3653 9854
rect 3579 9773 3590 9798
rect 3642 9773 3653 9798
rect 3579 9753 3653 9773
rect 3579 9701 3590 9753
rect 3642 9701 3653 9753
rect 3579 9663 3653 9701
rect 4095 9825 4169 9863
rect 4095 9773 4106 9825
rect 4158 9773 4169 9825
rect 4095 9753 4169 9773
rect 4095 9724 4106 9753
rect 4158 9724 4169 9753
rect 4095 9668 4104 9724
rect 4160 9668 4169 9724
rect 4095 9659 4169 9668
rect 4611 9854 4685 9863
rect 4611 9798 4620 9854
rect 4676 9798 4685 9854
rect 4611 9773 4622 9798
rect 4674 9773 4685 9798
rect 4611 9753 4685 9773
rect 4611 9701 4622 9753
rect 4674 9701 4685 9753
rect 4611 9659 4685 9701
rect 5621 9631 5667 9997
rect 9134 9688 9208 10400
rect 7335 9636 7351 9688
rect 7403 9636 7423 9688
rect 7475 9636 7609 9688
rect 7661 9636 7681 9688
rect 7733 9636 7867 9688
rect 7919 9636 7939 9688
rect 7991 9636 8125 9688
rect 8177 9636 8197 9688
rect 8249 9636 9208 9688
rect 3909 9628 3941 9631
rect 3907 9582 3941 9628
rect 3909 9579 3941 9582
rect 3993 9579 4013 9631
rect 4065 9579 4199 9631
rect 4251 9579 4271 9631
rect 4323 9579 5667 9631
rect 9134 9580 9208 9636
rect 2543 9474 3941 9526
rect 3993 9474 4013 9526
rect 4065 9474 4199 9526
rect 4251 9474 4271 9526
rect 4323 9474 4357 9526
rect 2543 9104 2589 9474
rect 3579 9407 3653 9445
rect 3579 9355 3590 9407
rect 3642 9355 3653 9407
rect 3579 9335 3653 9355
rect 3579 9306 3590 9335
rect 3642 9306 3653 9335
rect 3579 9250 3588 9306
rect 3644 9250 3653 9306
rect 3579 9241 3653 9250
rect 4095 9435 4169 9445
rect 4095 9379 4104 9435
rect 4160 9379 4169 9435
rect 4095 9355 4106 9379
rect 4158 9355 4169 9379
rect 4095 9335 4169 9355
rect 4095 9283 4106 9335
rect 4158 9283 4169 9335
rect 4095 9245 4169 9283
rect 4611 9407 4685 9445
rect 4611 9355 4622 9407
rect 4674 9355 4685 9407
rect 4611 9335 4685 9355
rect 4611 9306 4622 9335
rect 4674 9306 4685 9335
rect 4611 9250 4620 9306
rect 4676 9250 4685 9306
rect 4611 9241 4685 9250
rect 5621 9213 5667 9579
rect 7335 9528 7351 9580
rect 7403 9528 7423 9580
rect 7475 9528 7609 9580
rect 7661 9528 7681 9580
rect 7733 9528 7867 9580
rect 7919 9528 7939 9580
rect 7991 9528 8125 9580
rect 8177 9528 8197 9580
rect 8249 9528 9208 9580
rect 3391 9161 3425 9213
rect 3477 9161 3497 9213
rect 3549 9161 3683 9213
rect 3735 9161 3755 9213
rect 3807 9161 4457 9213
rect 4509 9161 4529 9213
rect 4581 9161 4715 9213
rect 4767 9161 4787 9213
rect 4839 9161 5667 9213
rect 2543 9052 3425 9104
rect 3477 9052 3497 9104
rect 3549 9052 3683 9104
rect 3735 9052 3755 9104
rect 3807 9052 4457 9104
rect 4509 9052 4529 9104
rect 4581 9052 4715 9104
rect 4767 9052 4787 9104
rect 4839 9052 4873 9104
rect 2543 8682 2589 9052
rect 3579 9014 3653 9023
rect 3579 8958 3588 9014
rect 3644 8958 3653 9014
rect 3579 8933 3590 8958
rect 3642 8933 3653 8958
rect 3579 8913 3653 8933
rect 3579 8861 3590 8913
rect 3642 8861 3653 8913
rect 3579 8823 3653 8861
rect 4095 8985 4169 9023
rect 4095 8933 4106 8985
rect 4158 8933 4169 8985
rect 4095 8913 4169 8933
rect 4095 8883 4106 8913
rect 4158 8883 4169 8913
rect 4095 8827 4104 8883
rect 4160 8827 4169 8883
rect 4095 8819 4169 8827
rect 4611 9014 4685 9023
rect 4611 8958 4620 9014
rect 4676 8958 4685 9014
rect 4611 8933 4622 8958
rect 4674 8933 4685 8958
rect 4611 8913 4685 8933
rect 4611 8861 4622 8913
rect 4674 8861 4685 8913
rect 4611 8823 4685 8861
rect 5621 8791 5667 9161
rect 9134 8816 9208 9528
rect 3907 8739 3941 8791
rect 3993 8739 4013 8791
rect 4065 8739 4199 8791
rect 4251 8739 4271 8791
rect 4323 8739 5667 8791
rect 7335 8764 7351 8816
rect 7403 8764 7423 8816
rect 7475 8764 7609 8816
rect 7661 8764 7681 8816
rect 7733 8764 7867 8816
rect 7919 8764 7939 8816
rect 7991 8764 8125 8816
rect 8177 8764 8197 8816
rect 8249 8764 9208 8816
rect 2543 8676 3941 8682
rect -5040 8630 3941 8676
rect 3993 8630 4013 8682
rect 4065 8630 4199 8682
rect 4251 8630 4271 8682
rect 4323 8630 4357 8682
rect 3579 8563 3653 8601
rect 3579 8511 3590 8563
rect 3642 8511 3653 8563
rect 3579 8491 3653 8511
rect 3579 8462 3590 8491
rect 3642 8462 3653 8491
rect 3579 8406 3588 8462
rect 3644 8406 3653 8462
rect 3579 8397 3653 8406
rect 4095 8592 4169 8601
rect 4095 8536 4104 8592
rect 4160 8536 4169 8592
rect 4095 8511 4106 8536
rect 4158 8511 4169 8536
rect 4095 8491 4169 8511
rect 4095 8439 4106 8491
rect 4158 8439 4169 8491
rect 4095 8401 4169 8439
rect 4611 8563 4685 8601
rect 4611 8511 4622 8563
rect 4674 8511 4685 8563
rect 4611 8491 4685 8511
rect 4611 8462 4622 8491
rect 4674 8462 4685 8491
rect 4611 8406 4620 8462
rect 4676 8406 4685 8462
rect 4611 8397 4685 8406
rect 2227 8374 2307 8383
rect 2227 8318 2239 8374
rect 2295 8318 2307 8374
rect 5621 8369 5667 8739
rect 9134 8708 9208 8764
rect 7335 8656 7351 8708
rect 7403 8656 7423 8708
rect 7475 8656 7609 8708
rect 7661 8656 7681 8708
rect 7733 8656 7867 8708
rect 7919 8656 7939 8708
rect 7991 8656 8125 8708
rect 8177 8656 8197 8708
rect 8249 8656 9208 8708
rect 2227 8307 2307 8318
rect 3649 8317 3683 8369
rect 3735 8317 3755 8369
rect 3807 8317 4457 8369
rect 4509 8317 4529 8369
rect 4581 8323 5667 8369
rect 4581 8317 5621 8323
rect 9134 8272 9208 8656
rect 7335 8220 7351 8272
rect 7403 8220 7423 8272
rect 7475 8220 7609 8272
rect 7661 8220 7681 8272
rect 7733 8220 7867 8272
rect 7919 8220 7939 8272
rect 7991 8220 8125 8272
rect 8177 8220 8197 8272
rect 8249 8220 9208 8272
rect -2942 8031 -2890 8163
rect -2942 7979 -834 8031
rect -782 7979 -762 8031
rect -710 7979 -576 8031
rect -524 7979 -504 8031
rect -452 7979 -318 8031
rect -266 7979 -246 8031
rect -194 7979 -60 8031
rect -8 7979 12 8031
rect 64 7979 198 8031
rect 250 7979 270 8031
rect 322 7979 456 8031
rect 508 7979 528 8031
rect 580 7979 596 8031
rect 3197 7985 3277 7994
rect -2942 7613 -2890 7979
rect -680 7941 -606 7950
rect -680 7885 -671 7941
rect -615 7885 -606 7941
rect -680 7860 -669 7885
rect -617 7860 -606 7885
rect -680 7840 -606 7860
rect -680 7788 -669 7840
rect -617 7788 -606 7840
rect -680 7750 -606 7788
rect -164 7941 -90 7950
rect -164 7885 -155 7941
rect -99 7885 -90 7941
rect -164 7860 -153 7885
rect -101 7860 -90 7885
rect -164 7840 -90 7860
rect -164 7788 -153 7840
rect -101 7788 -90 7840
rect -164 7750 -90 7788
rect 352 7941 426 7950
rect 352 7885 361 7941
rect 417 7885 426 7941
rect 3197 7929 3209 7985
rect 3265 7929 3277 7985
rect 9134 7960 9208 8220
rect 3197 7918 3277 7929
rect 352 7860 363 7885
rect 415 7860 426 7885
rect 352 7840 426 7860
rect 352 7788 363 7840
rect 415 7788 426 7840
rect 352 7750 426 7788
rect 1894 7682 6761 7742
rect -2942 7561 -1350 7613
rect -1298 7561 -1278 7613
rect -1226 7561 -1092 7613
rect -1040 7561 -1020 7613
rect -968 7561 -318 7613
rect -266 7561 -246 7613
rect -194 7561 -60 7613
rect -8 7561 12 7613
rect 64 7561 714 7613
rect 766 7561 786 7613
rect 838 7561 972 7613
rect 1024 7561 1044 7613
rect 1096 7561 1112 7613
rect -2942 7195 -2890 7561
rect -1196 7523 -1122 7532
rect -1196 7467 -1187 7523
rect -1131 7467 -1122 7523
rect -1196 7442 -1185 7467
rect -1133 7442 -1122 7467
rect -1196 7422 -1122 7442
rect -1196 7370 -1185 7422
rect -1133 7370 -1122 7422
rect -1196 7332 -1122 7370
rect -680 7494 -606 7532
rect -680 7442 -669 7494
rect -617 7442 -606 7494
rect -680 7422 -606 7442
rect -680 7397 -669 7422
rect -617 7397 -606 7422
rect -680 7341 -671 7397
rect -615 7341 -606 7397
rect -680 7332 -606 7341
rect -164 7523 -90 7532
rect -164 7467 -155 7523
rect -99 7467 -90 7523
rect -164 7442 -153 7467
rect -101 7442 -90 7467
rect -164 7422 -90 7442
rect -164 7370 -153 7422
rect -101 7370 -90 7422
rect -164 7332 -90 7370
rect 352 7494 426 7532
rect 352 7442 363 7494
rect 415 7442 426 7494
rect 352 7422 426 7442
rect 352 7397 363 7422
rect 415 7397 426 7422
rect 352 7341 361 7397
rect 417 7341 426 7397
rect 352 7332 426 7341
rect 868 7523 942 7532
rect 868 7467 877 7523
rect 933 7467 942 7523
rect 868 7442 879 7467
rect 931 7442 942 7467
rect 868 7422 942 7442
rect 868 7370 879 7422
rect 931 7370 942 7422
rect 868 7332 942 7370
rect 1894 7303 1940 7682
rect -1882 7251 -834 7303
rect -782 7251 -762 7303
rect -710 7251 -576 7303
rect -524 7251 -504 7303
rect -452 7251 198 7303
rect 250 7251 270 7303
rect 322 7251 456 7303
rect 508 7251 528 7303
rect 580 7251 1940 7303
rect -2942 7143 -1866 7195
rect -1814 7143 -1794 7195
rect -1742 7143 -1608 7195
rect -1556 7143 -1536 7195
rect -1484 7143 -834 7195
rect -782 7143 -762 7195
rect -710 7143 -576 7195
rect -524 7143 -504 7195
rect -452 7143 198 7195
rect 250 7143 270 7195
rect 322 7143 456 7195
rect 508 7143 528 7195
rect 580 7143 1112 7195
rect -2942 6777 -2890 7143
rect -1712 7105 -1638 7114
rect -1712 7049 -1703 7105
rect -1647 7049 -1638 7105
rect -1712 7024 -1701 7049
rect -1649 7024 -1638 7049
rect -1712 7004 -1638 7024
rect -1712 6952 -1701 7004
rect -1649 6952 -1638 7004
rect -1712 6914 -1638 6952
rect -1196 7076 -1122 7114
rect -1196 7024 -1185 7076
rect -1133 7024 -1122 7076
rect -1196 7004 -1122 7024
rect -1196 6979 -1185 7004
rect -1133 6979 -1122 7004
rect -1196 6923 -1187 6979
rect -1131 6923 -1122 6979
rect -1196 6914 -1122 6923
rect -680 7105 -606 7114
rect -680 7049 -671 7105
rect -615 7049 -606 7105
rect -680 7024 -669 7049
rect -617 7024 -606 7049
rect -680 7004 -606 7024
rect -680 6952 -669 7004
rect -617 6952 -606 7004
rect -680 6914 -606 6952
rect -164 7076 -90 7114
rect -164 7024 -153 7076
rect -101 7024 -90 7076
rect -164 7004 -90 7024
rect -164 6979 -153 7004
rect -101 6979 -90 7004
rect -164 6923 -155 6979
rect -99 6923 -90 6979
rect -164 6914 -90 6923
rect 352 7105 426 7114
rect 352 7049 361 7105
rect 417 7049 426 7105
rect 352 7024 363 7049
rect 415 7024 426 7049
rect 352 7004 426 7024
rect 352 6952 363 7004
rect 415 6952 426 7004
rect 352 6914 426 6952
rect 868 7076 942 7114
rect 868 7024 879 7076
rect 931 7024 942 7076
rect 868 7004 942 7024
rect 868 6979 879 7004
rect 931 6979 942 7004
rect 868 6923 877 6979
rect 933 6923 942 6979
rect 868 6914 942 6923
rect 1894 6885 1940 7251
rect -1882 6833 -1350 6885
rect -1298 6833 -1278 6885
rect -1226 6833 -1092 6885
rect -1040 6833 -1020 6885
rect -968 6833 -318 6885
rect -266 6833 -246 6885
rect -194 6833 -60 6885
rect -8 6833 12 6885
rect 64 6833 714 6885
rect 766 6833 786 6885
rect 838 6833 972 6885
rect 1024 6833 1044 6885
rect 1096 6833 1940 6885
rect -2942 6725 -1350 6777
rect -1298 6725 -1278 6777
rect -1226 6725 -1092 6777
rect -1040 6725 -1020 6777
rect -968 6725 -318 6777
rect -266 6725 -246 6777
rect -194 6725 -60 6777
rect -8 6725 12 6777
rect 64 6725 714 6777
rect 766 6725 786 6777
rect 838 6725 972 6777
rect 1024 6725 1044 6777
rect 1096 6725 1112 6777
rect -2942 6359 -2890 6725
rect -1712 6658 -1638 6696
rect -1712 6606 -1701 6658
rect -1649 6606 -1638 6658
rect -1712 6586 -1638 6606
rect -1712 6561 -1701 6586
rect -1649 6561 -1638 6586
rect -1712 6505 -1703 6561
rect -1647 6505 -1638 6561
rect -1712 6496 -1638 6505
rect -1196 6687 -1122 6696
rect -1196 6631 -1187 6687
rect -1131 6631 -1122 6687
rect -1196 6606 -1185 6631
rect -1133 6606 -1122 6631
rect -1196 6586 -1122 6606
rect -1196 6534 -1185 6586
rect -1133 6534 -1122 6586
rect -1196 6496 -1122 6534
rect -680 6658 -606 6696
rect -680 6606 -669 6658
rect -617 6606 -606 6658
rect -680 6586 -606 6606
rect -680 6561 -669 6586
rect -617 6561 -606 6586
rect -680 6505 -671 6561
rect -615 6505 -606 6561
rect -680 6496 -606 6505
rect -164 6687 -90 6696
rect -164 6631 -155 6687
rect -99 6631 -90 6687
rect -164 6606 -153 6631
rect -101 6606 -90 6631
rect -164 6586 -90 6606
rect -164 6534 -153 6586
rect -101 6534 -90 6586
rect -164 6496 -90 6534
rect 352 6658 426 6696
rect 352 6606 363 6658
rect 415 6606 426 6658
rect 352 6586 426 6606
rect 352 6561 363 6586
rect 415 6561 426 6586
rect 352 6505 361 6561
rect 417 6505 426 6561
rect 352 6496 426 6505
rect 868 6687 942 6696
rect 868 6631 877 6687
rect 933 6631 942 6687
rect 868 6606 879 6631
rect 931 6606 942 6631
rect 868 6586 942 6606
rect 868 6534 879 6586
rect 931 6534 942 6586
rect 868 6496 942 6534
rect 1894 6467 1940 6833
rect -1882 6415 -1866 6467
rect -1814 6415 -1794 6467
rect -1742 6415 -1608 6467
rect -1556 6415 -1536 6467
rect -1484 6415 -834 6467
rect -782 6415 -762 6467
rect -710 6415 -576 6467
rect -524 6415 -504 6467
rect -452 6415 198 6467
rect 250 6415 270 6467
rect 322 6415 456 6467
rect 508 6415 528 6467
rect 580 6415 1940 6467
rect -2942 6307 -1866 6359
rect -1814 6307 -1794 6359
rect -1742 6307 -1608 6359
rect -1556 6307 -1536 6359
rect -1484 6307 -834 6359
rect -782 6307 -762 6359
rect -710 6307 -576 6359
rect -524 6307 -504 6359
rect -452 6307 198 6359
rect 250 6307 270 6359
rect 322 6307 456 6359
rect 508 6307 528 6359
rect 580 6307 1112 6359
rect -2942 5941 -2890 6307
rect -1712 6269 -1638 6278
rect -1712 6213 -1703 6269
rect -1647 6213 -1638 6269
rect -1712 6188 -1701 6213
rect -1649 6188 -1638 6213
rect -1712 6168 -1638 6188
rect -1712 6116 -1701 6168
rect -1649 6116 -1638 6168
rect -1712 6078 -1638 6116
rect -1196 6240 -1122 6278
rect -1196 6188 -1185 6240
rect -1133 6188 -1122 6240
rect -1196 6168 -1122 6188
rect -1196 6143 -1185 6168
rect -1133 6143 -1122 6168
rect -1196 6087 -1187 6143
rect -1131 6087 -1122 6143
rect -1196 6078 -1122 6087
rect -680 6269 -606 6278
rect -680 6213 -671 6269
rect -615 6213 -606 6269
rect -680 6188 -669 6213
rect -617 6188 -606 6213
rect -680 6168 -606 6188
rect -680 6116 -669 6168
rect -617 6116 -606 6168
rect -680 6078 -606 6116
rect -164 6240 -90 6278
rect -164 6188 -153 6240
rect -101 6188 -90 6240
rect -164 6168 -90 6188
rect -164 6143 -153 6168
rect -101 6143 -90 6168
rect -164 6087 -155 6143
rect -99 6087 -90 6143
rect -164 6078 -90 6087
rect 352 6269 426 6278
rect 352 6213 361 6269
rect 417 6213 426 6269
rect 352 6188 363 6213
rect 415 6188 426 6213
rect 352 6168 426 6188
rect 352 6116 363 6168
rect 415 6116 426 6168
rect 352 6078 426 6116
rect 868 6240 942 6278
rect 868 6188 879 6240
rect 931 6188 942 6240
rect 868 6168 942 6188
rect 868 6143 879 6168
rect 931 6143 942 6168
rect 868 6087 877 6143
rect 933 6087 942 6143
rect 868 6078 942 6087
rect 1894 6049 1940 6415
rect -1882 5997 -1350 6049
rect -1298 5997 -1278 6049
rect -1226 5997 -1092 6049
rect -1040 5997 -1020 6049
rect -968 5997 -318 6049
rect -266 5997 -246 6049
rect -194 5997 -60 6049
rect -8 5997 12 6049
rect 64 5997 714 6049
rect 766 5997 786 6049
rect 838 5997 972 6049
rect 1024 5997 1044 6049
rect 1096 5997 1940 6049
rect -2942 5889 -1350 5941
rect -1298 5889 -1278 5941
rect -1226 5889 -1092 5941
rect -1040 5889 -1020 5941
rect -968 5889 -318 5941
rect -266 5889 -246 5941
rect -194 5889 -60 5941
rect -8 5889 12 5941
rect 64 5889 714 5941
rect 766 5889 786 5941
rect 838 5889 972 5941
rect 1024 5889 1044 5941
rect 1096 5889 1112 5941
rect -2942 5523 -2890 5889
rect -1712 5822 -1638 5860
rect -1712 5770 -1701 5822
rect -1649 5770 -1638 5822
rect -1712 5750 -1638 5770
rect -1712 5725 -1701 5750
rect -1649 5725 -1638 5750
rect -1712 5669 -1703 5725
rect -1647 5669 -1638 5725
rect -1712 5660 -1638 5669
rect -1196 5851 -1122 5860
rect -1196 5795 -1187 5851
rect -1131 5795 -1122 5851
rect -1196 5770 -1185 5795
rect -1133 5770 -1122 5795
rect -1196 5750 -1122 5770
rect -1196 5698 -1185 5750
rect -1133 5698 -1122 5750
rect -1196 5660 -1122 5698
rect -680 5822 -606 5860
rect -680 5770 -669 5822
rect -617 5770 -606 5822
rect -680 5750 -606 5770
rect -680 5725 -669 5750
rect -617 5725 -606 5750
rect -680 5669 -671 5725
rect -615 5669 -606 5725
rect -680 5660 -606 5669
rect -164 5851 -90 5860
rect -164 5795 -155 5851
rect -99 5795 -90 5851
rect -164 5770 -153 5795
rect -101 5770 -90 5795
rect -164 5750 -90 5770
rect -164 5698 -153 5750
rect -101 5698 -90 5750
rect -164 5660 -90 5698
rect 352 5822 426 5860
rect 352 5770 363 5822
rect 415 5770 426 5822
rect 352 5750 426 5770
rect 352 5725 363 5750
rect 415 5725 426 5750
rect 352 5669 361 5725
rect 417 5669 426 5725
rect 352 5660 426 5669
rect 868 5851 942 5860
rect 868 5795 877 5851
rect 933 5795 942 5851
rect 868 5770 879 5795
rect 931 5770 942 5795
rect 868 5750 942 5770
rect 868 5698 879 5750
rect 931 5698 942 5750
rect 868 5660 942 5698
rect 1894 5631 1940 5997
rect -1882 5579 -1866 5631
rect -1814 5579 -1794 5631
rect -1742 5579 -1608 5631
rect -1556 5579 -1536 5631
rect -1484 5579 -834 5631
rect -782 5579 -762 5631
rect -710 5579 -576 5631
rect -524 5579 -504 5631
rect -452 5579 198 5631
rect 250 5579 270 5631
rect 322 5579 456 5631
rect 508 5579 528 5631
rect 580 5579 1940 5631
rect -2942 5471 -1866 5523
rect -1814 5471 -1794 5523
rect -1742 5471 -1608 5523
rect -1556 5471 -1536 5523
rect -1484 5471 -834 5523
rect -782 5471 -762 5523
rect -710 5471 -576 5523
rect -524 5471 -504 5523
rect -452 5471 198 5523
rect 250 5471 270 5523
rect 322 5471 456 5523
rect 508 5471 528 5523
rect 580 5471 1112 5523
rect -2942 5105 -2890 5471
rect -1712 5433 -1638 5442
rect -1712 5377 -1703 5433
rect -1647 5377 -1638 5433
rect -1712 5352 -1701 5377
rect -1649 5352 -1638 5377
rect -1712 5332 -1638 5352
rect -1712 5280 -1701 5332
rect -1649 5280 -1638 5332
rect -1712 5242 -1638 5280
rect -1196 5404 -1122 5442
rect -1196 5352 -1185 5404
rect -1133 5352 -1122 5404
rect -1196 5332 -1122 5352
rect -1196 5307 -1185 5332
rect -1133 5307 -1122 5332
rect -1196 5251 -1187 5307
rect -1131 5251 -1122 5307
rect -1196 5242 -1122 5251
rect -680 5433 -606 5442
rect -680 5377 -671 5433
rect -615 5377 -606 5433
rect -680 5352 -669 5377
rect -617 5352 -606 5377
rect -680 5332 -606 5352
rect -680 5280 -669 5332
rect -617 5280 -606 5332
rect -680 5242 -606 5280
rect -164 5404 -90 5442
rect -164 5352 -153 5404
rect -101 5352 -90 5404
rect -164 5332 -90 5352
rect -164 5307 -153 5332
rect -101 5307 -90 5332
rect -164 5251 -155 5307
rect -99 5251 -90 5307
rect -164 5242 -90 5251
rect 352 5433 426 5442
rect 352 5377 361 5433
rect 417 5377 426 5433
rect 352 5352 363 5377
rect 415 5352 426 5377
rect 352 5332 426 5352
rect 352 5280 363 5332
rect 415 5280 426 5332
rect 352 5242 426 5280
rect 868 5404 942 5442
rect 868 5352 879 5404
rect 931 5352 942 5404
rect 868 5332 942 5352
rect 868 5307 879 5332
rect 931 5307 942 5332
rect 868 5251 877 5307
rect 933 5251 942 5307
rect 868 5242 942 5251
rect 1894 5213 1940 5579
rect -1882 5161 -1350 5213
rect -1298 5161 -1278 5213
rect -1226 5161 -1092 5213
rect -1040 5161 -1020 5213
rect -968 5161 -318 5213
rect -266 5161 -246 5213
rect -194 5161 -60 5213
rect -8 5161 12 5213
rect 64 5161 714 5213
rect 766 5161 786 5213
rect 838 5161 972 5213
rect 1024 5161 1044 5213
rect 1096 5161 1940 5213
rect -2942 5053 -1350 5105
rect -1298 5053 -1278 5105
rect -1226 5053 -1092 5105
rect -1040 5053 -1020 5105
rect -968 5053 -318 5105
rect -266 5053 -246 5105
rect -194 5053 -60 5105
rect -8 5053 12 5105
rect 64 5053 714 5105
rect 766 5053 786 5105
rect 838 5053 972 5105
rect 1024 5053 1044 5105
rect 1096 5053 1112 5105
rect -2942 4687 -2890 5053
rect -1712 4986 -1638 5024
rect -1712 4934 -1701 4986
rect -1649 4934 -1638 4986
rect -1712 4914 -1638 4934
rect -1712 4889 -1701 4914
rect -1649 4889 -1638 4914
rect -1712 4833 -1703 4889
rect -1647 4833 -1638 4889
rect -1712 4824 -1638 4833
rect -1196 5015 -1122 5024
rect -1196 4959 -1187 5015
rect -1131 4959 -1122 5015
rect -1196 4934 -1185 4959
rect -1133 4934 -1122 4959
rect -1196 4914 -1122 4934
rect -1196 4862 -1185 4914
rect -1133 4862 -1122 4914
rect -1196 4824 -1122 4862
rect -680 4986 -606 5024
rect -680 4934 -669 4986
rect -617 4934 -606 4986
rect -680 4914 -606 4934
rect -680 4889 -669 4914
rect -617 4889 -606 4914
rect -680 4833 -671 4889
rect -615 4833 -606 4889
rect -680 4824 -606 4833
rect -164 5015 -90 5024
rect -164 4959 -155 5015
rect -99 4959 -90 5015
rect -164 4934 -153 4959
rect -101 4934 -90 4959
rect -164 4914 -90 4934
rect -164 4862 -153 4914
rect -101 4862 -90 4914
rect -164 4824 -90 4862
rect 352 4986 426 5024
rect 352 4934 363 4986
rect 415 4934 426 4986
rect 352 4914 426 4934
rect 352 4889 363 4914
rect 415 4889 426 4914
rect 352 4833 361 4889
rect 417 4833 426 4889
rect 352 4824 426 4833
rect 868 5015 942 5024
rect 868 4959 877 5015
rect 933 4959 942 5015
rect 868 4934 879 4959
rect 931 4934 942 4959
rect 868 4914 942 4934
rect 868 4862 879 4914
rect 931 4862 942 4914
rect 868 4824 942 4862
rect 1894 4795 1940 5161
rect -1882 4743 -1866 4795
rect -1814 4743 -1794 4795
rect -1742 4743 -1608 4795
rect -1556 4743 -1536 4795
rect -1484 4743 -834 4795
rect -782 4743 -762 4795
rect -710 4743 -576 4795
rect -524 4743 -504 4795
rect -452 4743 198 4795
rect 250 4743 270 4795
rect 322 4743 456 4795
rect 508 4743 528 4795
rect 580 4743 1940 4795
rect -2942 4635 -1866 4687
rect -1814 4635 -1794 4687
rect -1742 4635 -1608 4687
rect -1556 4635 -1536 4687
rect -1484 4635 -834 4687
rect -782 4635 -762 4687
rect -710 4635 -576 4687
rect -524 4635 -504 4687
rect -452 4635 198 4687
rect 250 4635 270 4687
rect 322 4635 456 4687
rect 508 4635 528 4687
rect 580 4635 1112 4687
rect -2942 4269 -2890 4635
rect -1712 4597 -1638 4606
rect -1712 4541 -1703 4597
rect -1647 4541 -1638 4597
rect -1712 4516 -1701 4541
rect -1649 4516 -1638 4541
rect -1712 4496 -1638 4516
rect -1712 4444 -1701 4496
rect -1649 4444 -1638 4496
rect -1712 4406 -1638 4444
rect -1196 4568 -1122 4606
rect -1196 4516 -1185 4568
rect -1133 4516 -1122 4568
rect -1196 4496 -1122 4516
rect -1196 4471 -1185 4496
rect -1133 4471 -1122 4496
rect -1196 4415 -1187 4471
rect -1131 4415 -1122 4471
rect -1196 4406 -1122 4415
rect -680 4597 -606 4606
rect -680 4541 -671 4597
rect -615 4541 -606 4597
rect -680 4516 -669 4541
rect -617 4516 -606 4541
rect -680 4496 -606 4516
rect -680 4444 -669 4496
rect -617 4444 -606 4496
rect -680 4406 -606 4444
rect -164 4568 -90 4606
rect -164 4516 -153 4568
rect -101 4516 -90 4568
rect -164 4496 -90 4516
rect -164 4471 -153 4496
rect -101 4471 -90 4496
rect -164 4415 -155 4471
rect -99 4415 -90 4471
rect -164 4406 -90 4415
rect 352 4597 426 4606
rect 352 4541 361 4597
rect 417 4541 426 4597
rect 352 4516 363 4541
rect 415 4516 426 4541
rect 352 4496 426 4516
rect 352 4444 363 4496
rect 415 4444 426 4496
rect 352 4406 426 4444
rect 1894 4377 1940 4743
rect -1882 4325 -1350 4377
rect -1298 4325 -1278 4377
rect -1226 4325 -1092 4377
rect -1040 4325 -1020 4377
rect -968 4325 -318 4377
rect -266 4325 -246 4377
rect -194 4325 -60 4377
rect -8 4325 12 4377
rect 64 4325 1940 4377
rect -2942 4217 -1350 4269
rect -1298 4217 -1278 4269
rect -1226 4217 -1092 4269
rect -1040 4217 -1020 4269
rect -968 4217 -834 4269
rect -782 4217 -762 4269
rect -710 4217 -576 4269
rect -524 4217 -504 4269
rect -452 4217 -318 4269
rect -266 4217 -246 4269
rect -194 4217 -60 4269
rect -8 4217 12 4269
rect 64 4217 1112 4269
rect -2942 3668 -2890 4217
rect 1894 4204 1940 4325
rect 2891 7392 2943 7525
rect 2891 7340 3964 7392
rect 4016 7340 4036 7392
rect 4088 7340 4222 7392
rect 4274 7340 4294 7392
rect 4346 7340 4480 7392
rect 4532 7340 4552 7392
rect 4604 7340 4738 7392
rect 4790 7340 4810 7392
rect 4862 7340 4996 7392
rect 5048 7340 5068 7392
rect 5120 7340 5254 7392
rect 5306 7340 5326 7392
rect 5378 7340 5512 7392
rect 5564 7340 5584 7392
rect 5636 7340 5770 7392
rect 5822 7340 5842 7392
rect 5894 7340 5910 7392
rect 2891 6974 2943 7340
rect 4118 7302 4192 7311
rect 4118 7246 4127 7302
rect 4183 7246 4192 7302
rect 4118 7221 4129 7246
rect 4181 7221 4192 7246
rect 4118 7201 4192 7221
rect 4118 7149 4129 7201
rect 4181 7149 4192 7201
rect 4118 7111 4192 7149
rect 4634 7302 4708 7311
rect 4634 7246 4643 7302
rect 4699 7246 4708 7302
rect 4634 7221 4645 7246
rect 4697 7221 4708 7246
rect 4634 7201 4708 7221
rect 4634 7149 4645 7201
rect 4697 7149 4708 7201
rect 4634 7111 4708 7149
rect 5150 7302 5224 7311
rect 5150 7246 5159 7302
rect 5215 7246 5224 7302
rect 5150 7221 5161 7246
rect 5213 7221 5224 7246
rect 5150 7201 5224 7221
rect 5150 7149 5161 7201
rect 5213 7149 5224 7201
rect 5150 7111 5224 7149
rect 5666 7302 5740 7311
rect 5666 7246 5675 7302
rect 5731 7246 5740 7302
rect 5666 7221 5677 7246
rect 5729 7221 5740 7246
rect 5666 7201 5740 7221
rect 5666 7149 5677 7201
rect 5729 7149 5740 7201
rect 5666 7111 5740 7149
rect 2891 6922 3964 6974
rect 4016 6922 4036 6974
rect 4088 6922 4222 6974
rect 4274 6922 4294 6974
rect 4346 6922 4996 6974
rect 5048 6922 5068 6974
rect 5120 6922 5254 6974
rect 5306 6922 5326 6974
rect 5378 6922 5910 6974
rect 2891 6556 2943 6922
rect 4118 6884 4192 6893
rect 4118 6828 4127 6884
rect 4183 6828 4192 6884
rect 4118 6803 4129 6828
rect 4181 6803 4192 6828
rect 4118 6783 4192 6803
rect 4118 6731 4129 6783
rect 4181 6731 4192 6783
rect 4118 6693 4192 6731
rect 4634 6855 4708 6893
rect 4634 6803 4645 6855
rect 4697 6803 4708 6855
rect 4634 6783 4708 6803
rect 4634 6758 4645 6783
rect 4697 6758 4708 6783
rect 4634 6702 4643 6758
rect 4699 6702 4708 6758
rect 4634 6693 4708 6702
rect 5150 6884 5224 6893
rect 5150 6828 5159 6884
rect 5215 6828 5224 6884
rect 5150 6803 5161 6828
rect 5213 6803 5224 6828
rect 5150 6783 5224 6803
rect 5150 6731 5161 6783
rect 5213 6731 5224 6783
rect 5150 6693 5224 6731
rect 5666 6855 5740 6893
rect 5666 6803 5677 6855
rect 5729 6803 5740 6855
rect 5666 6783 5740 6803
rect 5666 6758 5677 6783
rect 5729 6758 5740 6783
rect 5666 6702 5675 6758
rect 5731 6702 5740 6758
rect 5666 6693 5740 6702
rect 6701 6664 6761 7682
rect 7774 7283 12290 7343
rect 7774 6981 7834 7283
rect 7630 6929 8700 6981
rect 8752 6929 8772 6981
rect 8824 6929 8958 6981
rect 9010 6929 9030 6981
rect 9082 6929 9216 6981
rect 9268 6929 9288 6981
rect 9340 6929 9474 6981
rect 9526 6929 9546 6981
rect 9598 6929 9614 6981
rect 7630 6664 7676 6929
rect 8596 6810 8607 6862
rect 8659 6810 9123 6862
rect 9175 6810 9639 6862
rect 9691 6810 9704 6862
rect 3948 6612 4480 6664
rect 4532 6612 4552 6664
rect 4604 6612 4738 6664
rect 4790 6612 4810 6664
rect 4862 6612 5512 6664
rect 5564 6612 5584 6664
rect 5636 6612 5770 6664
rect 5822 6612 5842 6664
rect 5894 6612 7676 6664
rect 6918 6604 7676 6612
rect 2891 6504 4480 6556
rect 4532 6504 4552 6556
rect 4604 6504 4738 6556
rect 4790 6504 4810 6556
rect 4862 6504 5512 6556
rect 5564 6504 5584 6556
rect 5636 6504 5770 6556
rect 5822 6504 5842 6556
rect 5894 6504 5910 6556
rect 2891 6138 2943 6504
rect 4118 6437 4192 6475
rect 4118 6385 4129 6437
rect 4181 6385 4192 6437
rect 4118 6365 4192 6385
rect 4118 6340 4129 6365
rect 4181 6340 4192 6365
rect 4118 6284 4127 6340
rect 4183 6284 4192 6340
rect 4118 6275 4192 6284
rect 4634 6466 4708 6475
rect 4634 6410 4643 6466
rect 4699 6410 4708 6466
rect 4634 6385 4645 6410
rect 4697 6385 4708 6410
rect 4634 6365 4708 6385
rect 4634 6313 4645 6365
rect 4697 6313 4708 6365
rect 4634 6275 4708 6313
rect 5150 6437 5224 6475
rect 5150 6385 5161 6437
rect 5213 6385 5224 6437
rect 5150 6365 5224 6385
rect 5150 6340 5161 6365
rect 5213 6340 5224 6365
rect 5150 6284 5159 6340
rect 5215 6284 5224 6340
rect 5150 6275 5224 6284
rect 5666 6466 5740 6475
rect 5666 6410 5675 6466
rect 5731 6410 5740 6466
rect 5666 6385 5677 6410
rect 5729 6385 5740 6410
rect 5666 6365 5740 6385
rect 5666 6313 5677 6365
rect 5729 6313 5740 6365
rect 5666 6275 5740 6313
rect 6918 6246 6964 6604
rect 3948 6194 3964 6246
rect 4016 6194 4036 6246
rect 4088 6194 4222 6246
rect 4274 6194 4294 6246
rect 4346 6194 4996 6246
rect 5048 6194 5068 6246
rect 5120 6194 5254 6246
rect 5306 6194 5326 6246
rect 5378 6194 6964 6246
rect 2891 6086 3964 6138
rect 4016 6086 4036 6138
rect 4088 6086 4222 6138
rect 4274 6086 4294 6138
rect 4346 6086 4996 6138
rect 5048 6086 5068 6138
rect 5120 6086 5254 6138
rect 5306 6086 5326 6138
rect 5378 6086 5910 6138
rect 2891 5720 2943 6086
rect 4118 6048 4192 6057
rect 4118 5992 4127 6048
rect 4183 5992 4192 6048
rect 4118 5967 4129 5992
rect 4181 5967 4192 5992
rect 4118 5947 4192 5967
rect 4118 5895 4129 5947
rect 4181 5895 4192 5947
rect 4118 5857 4192 5895
rect 4634 6019 4708 6057
rect 4634 5967 4645 6019
rect 4697 5967 4708 6019
rect 4634 5947 4708 5967
rect 4634 5922 4645 5947
rect 4697 5922 4708 5947
rect 4634 5866 4643 5922
rect 4699 5866 4708 5922
rect 4634 5857 4708 5866
rect 5150 6048 5224 6057
rect 5150 5992 5159 6048
rect 5215 5992 5224 6048
rect 5150 5967 5161 5992
rect 5213 5967 5224 5992
rect 5150 5947 5224 5967
rect 5150 5895 5161 5947
rect 5213 5895 5224 5947
rect 5150 5857 5224 5895
rect 5666 6019 5740 6057
rect 5666 5967 5677 6019
rect 5729 5967 5740 6019
rect 5666 5947 5740 5967
rect 5666 5922 5677 5947
rect 5729 5922 5740 5947
rect 5666 5866 5675 5922
rect 5731 5866 5740 5922
rect 5666 5857 5740 5866
rect 6918 5828 6964 6194
rect 3948 5776 4480 5828
rect 4532 5776 4552 5828
rect 4604 5776 4738 5828
rect 4790 5776 4810 5828
rect 4862 5776 5512 5828
rect 5564 5776 5584 5828
rect 5636 5776 5770 5828
rect 5822 5776 5842 5828
rect 5894 5776 6964 5828
rect 2891 5668 4480 5720
rect 4532 5668 4552 5720
rect 4604 5668 4738 5720
rect 4790 5668 4810 5720
rect 4862 5668 5512 5720
rect 5564 5668 5584 5720
rect 5636 5668 5770 5720
rect 5822 5668 5842 5720
rect 5894 5668 5910 5720
rect 2891 5302 2943 5668
rect 4118 5601 4192 5639
rect 4118 5549 4129 5601
rect 4181 5549 4192 5601
rect 4118 5529 4192 5549
rect 4118 5504 4129 5529
rect 4181 5504 4192 5529
rect 4118 5448 4127 5504
rect 4183 5448 4192 5504
rect 4118 5439 4192 5448
rect 4634 5630 4708 5639
rect 4634 5574 4643 5630
rect 4699 5574 4708 5630
rect 4634 5549 4645 5574
rect 4697 5549 4708 5574
rect 4634 5529 4708 5549
rect 4634 5477 4645 5529
rect 4697 5477 4708 5529
rect 4634 5439 4708 5477
rect 5150 5601 5224 5639
rect 5150 5549 5161 5601
rect 5213 5549 5224 5601
rect 5150 5529 5224 5549
rect 5150 5504 5161 5529
rect 5213 5504 5224 5529
rect 5150 5448 5159 5504
rect 5215 5448 5224 5504
rect 5150 5439 5224 5448
rect 5666 5630 5740 5639
rect 5666 5574 5675 5630
rect 5731 5574 5740 5630
rect 5666 5549 5677 5574
rect 5729 5549 5740 5574
rect 5666 5529 5740 5549
rect 5666 5477 5677 5529
rect 5729 5477 5740 5529
rect 5666 5439 5740 5477
rect 6918 5410 6964 5776
rect 3948 5358 3964 5410
rect 4016 5358 4036 5410
rect 4088 5358 4222 5410
rect 4274 5358 4294 5410
rect 4346 5358 4996 5410
rect 5048 5358 5068 5410
rect 5120 5358 5254 5410
rect 5306 5358 5326 5410
rect 5378 5358 6964 5410
rect 2891 5250 3964 5302
rect 4016 5250 4036 5302
rect 4088 5250 4222 5302
rect 4274 5250 4294 5302
rect 4346 5250 4996 5302
rect 5048 5250 5068 5302
rect 5120 5250 5254 5302
rect 5306 5250 5326 5302
rect 5378 5250 5910 5302
rect 2891 4884 2943 5250
rect 4118 5212 4192 5221
rect 4118 5156 4127 5212
rect 4183 5156 4192 5212
rect 4118 5131 4129 5156
rect 4181 5131 4192 5156
rect 4118 5111 4192 5131
rect 4118 5059 4129 5111
rect 4181 5059 4192 5111
rect 4118 5021 4192 5059
rect 4634 5183 4708 5221
rect 4634 5131 4645 5183
rect 4697 5131 4708 5183
rect 4634 5111 4708 5131
rect 4634 5086 4645 5111
rect 4697 5086 4708 5111
rect 4634 5030 4643 5086
rect 4699 5030 4708 5086
rect 4634 5021 4708 5030
rect 5150 5212 5224 5221
rect 5150 5156 5159 5212
rect 5215 5156 5224 5212
rect 5150 5131 5161 5156
rect 5213 5131 5224 5156
rect 5150 5111 5224 5131
rect 5150 5059 5161 5111
rect 5213 5059 5224 5111
rect 5150 5021 5224 5059
rect 5666 5183 5740 5221
rect 5666 5131 5677 5183
rect 5729 5131 5740 5183
rect 5666 5111 5740 5131
rect 5666 5086 5677 5111
rect 5729 5086 5740 5111
rect 5666 5030 5675 5086
rect 5731 5030 5740 5086
rect 5666 5021 5740 5030
rect 6918 4992 6964 5358
rect 3948 4940 4480 4992
rect 4532 4940 4552 4992
rect 4604 4940 4738 4992
rect 4790 4940 4810 4992
rect 4862 4940 5512 4992
rect 5564 4940 5584 4992
rect 5636 4940 5770 4992
rect 5822 4940 5842 4992
rect 5894 4940 6964 4992
rect 2891 4832 4480 4884
rect 4532 4832 4552 4884
rect 4604 4832 4738 4884
rect 4790 4832 4810 4884
rect 4862 4832 5512 4884
rect 5564 4832 5584 4884
rect 5636 4832 5770 4884
rect 5822 4832 5842 4884
rect 5894 4832 5910 4884
rect 2891 4466 2943 4832
rect 4118 4765 4192 4803
rect 4118 4713 4129 4765
rect 4181 4713 4192 4765
rect 4118 4693 4192 4713
rect 4118 4668 4129 4693
rect 4181 4668 4192 4693
rect 4118 4612 4127 4668
rect 4183 4612 4192 4668
rect 4118 4603 4192 4612
rect 4634 4794 4708 4803
rect 4634 4738 4643 4794
rect 4699 4738 4708 4794
rect 4634 4713 4645 4738
rect 4697 4713 4708 4738
rect 4634 4693 4708 4713
rect 4634 4641 4645 4693
rect 4697 4641 4708 4693
rect 4634 4603 4708 4641
rect 5150 4765 5224 4803
rect 5150 4713 5161 4765
rect 5213 4713 5224 4765
rect 5150 4693 5224 4713
rect 5150 4668 5161 4693
rect 5213 4668 5224 4693
rect 5150 4612 5159 4668
rect 5215 4612 5224 4668
rect 5150 4603 5224 4612
rect 5666 4794 5740 4803
rect 5666 4738 5675 4794
rect 5731 4738 5740 4794
rect 5666 4713 5677 4738
rect 5729 4713 5740 4738
rect 5666 4693 5740 4713
rect 5666 4641 5677 4693
rect 5729 4641 5740 4693
rect 5666 4603 5740 4641
rect 6918 4574 6964 4940
rect 3948 4522 3964 4574
rect 4016 4522 4036 4574
rect 4088 4522 4222 4574
rect 4274 4522 4294 4574
rect 4346 4522 4996 4574
rect 5048 4522 5068 4574
rect 5120 4522 5254 4574
rect 5306 4522 5326 4574
rect 5378 4522 6964 4574
rect 2891 4414 3964 4466
rect 4016 4414 4036 4466
rect 4088 4414 4222 4466
rect 4274 4414 4294 4466
rect 4346 4414 4480 4466
rect 4532 4414 4552 4466
rect 4604 4414 4738 4466
rect 4790 4414 4810 4466
rect 4862 4414 4996 4466
rect 5048 4414 5068 4466
rect 5120 4414 5254 4466
rect 5306 4414 5326 4466
rect 5378 4414 5512 4466
rect 5564 4414 5584 4466
rect 5636 4414 5770 4466
rect 5822 4414 5842 4466
rect 5894 4414 5910 4466
rect -1196 4179 -1122 4188
rect -1196 4123 -1187 4179
rect -1131 4123 -1122 4179
rect -1196 4098 -1185 4123
rect -1133 4098 -1122 4123
rect -1196 4078 -1122 4098
rect -1196 4026 -1185 4078
rect -1133 4026 -1122 4078
rect -1196 3988 -1122 4026
rect -680 4179 -606 4188
rect -680 4123 -671 4179
rect -615 4123 -606 4179
rect -680 4098 -669 4123
rect -617 4098 -606 4123
rect -680 4078 -606 4098
rect -680 4026 -669 4078
rect -617 4026 -606 4078
rect -680 3988 -606 4026
rect -164 4179 -90 4188
rect -164 4123 -155 4179
rect -99 4123 -90 4179
rect -164 4098 -153 4123
rect -101 4098 -90 4123
rect -164 4078 -90 4098
rect -164 4026 -153 4078
rect -101 4026 -90 4078
rect -164 3988 -90 4026
rect 1381 4053 1461 4063
rect 1381 3997 1393 4053
rect 1449 3997 1461 4053
rect 1381 3987 1461 3997
rect 1495 4053 1575 4063
rect 1495 3997 1507 4053
rect 1563 3997 1575 4053
rect 1495 3987 1575 3997
rect 2891 3672 2943 4414
rect 6918 4407 6964 4522
rect 7630 6563 7676 6604
rect 7630 6511 8700 6563
rect 8752 6511 8772 6563
rect 8824 6511 8958 6563
rect 9010 6511 9030 6563
rect 9082 6511 9216 6563
rect 9268 6511 9288 6563
rect 9340 6511 9474 6563
rect 9526 6511 9546 6563
rect 9598 6511 9614 6563
rect 7630 6145 7676 6511
rect 7630 6093 8700 6145
rect 8752 6093 8772 6145
rect 8824 6093 8958 6145
rect 9010 6093 9030 6145
rect 9082 6093 9216 6145
rect 9268 6093 9288 6145
rect 9340 6093 9474 6145
rect 9526 6093 9546 6145
rect 9598 6093 9614 6145
rect 7630 5309 7676 6093
rect 8596 5675 8700 5727
rect 8752 5675 8772 5727
rect 8824 5675 8958 5727
rect 9010 5675 9030 5727
rect 9082 5675 9216 5727
rect 9268 5675 9288 5727
rect 9340 5675 9474 5727
rect 9526 5675 9546 5727
rect 9598 5675 12325 5727
rect 8596 5608 8670 5675
rect 8596 5556 8607 5608
rect 8659 5556 8670 5608
rect 8596 5536 8670 5556
rect 8596 5484 8607 5536
rect 8659 5484 8670 5536
rect 8596 5446 8670 5484
rect 9112 5608 9186 5675
rect 9112 5556 9123 5608
rect 9175 5556 9186 5608
rect 9112 5536 9186 5556
rect 9112 5484 9123 5536
rect 9175 5484 9186 5536
rect 9112 5446 9186 5484
rect 9628 5608 9702 5675
rect 9628 5556 9639 5608
rect 9691 5556 9702 5608
rect 9628 5536 9702 5556
rect 9628 5484 9639 5536
rect 9691 5484 9702 5536
rect 9628 5446 9702 5484
rect 7630 5257 8700 5309
rect 8752 5257 8772 5309
rect 8824 5257 8958 5309
rect 9010 5257 9030 5309
rect 9082 5257 9216 5309
rect 9268 5257 9288 5309
rect 9340 5257 9474 5309
rect 9526 5257 9546 5309
rect 9598 5257 9614 5309
rect 7630 4891 7676 5257
rect 7630 4839 8700 4891
rect 8752 4839 8772 4891
rect 8824 4839 8958 4891
rect 9010 4839 9030 4891
rect 9082 4839 9216 4891
rect 9268 4839 9288 4891
rect 9340 4839 9474 4891
rect 9526 4839 9546 4891
rect 9598 4839 9614 4891
rect 7630 4473 7676 4839
rect 7630 4421 8700 4473
rect 8752 4421 8772 4473
rect 8824 4421 8958 4473
rect 9010 4421 9030 4473
rect 9082 4421 9216 4473
rect 9268 4421 9288 4473
rect 9340 4421 9474 4473
rect 9526 4421 9546 4473
rect 9598 4421 9614 4473
rect 4118 4376 4192 4385
rect 4118 4320 4127 4376
rect 4183 4320 4192 4376
rect 4118 4295 4129 4320
rect 4181 4295 4192 4320
rect 4118 4275 4192 4295
rect 4118 4223 4129 4275
rect 4181 4223 4192 4275
rect 4118 4185 4192 4223
rect 4634 4376 4708 4385
rect 4634 4320 4643 4376
rect 4699 4320 4708 4376
rect 4634 4295 4645 4320
rect 4697 4295 4708 4320
rect 4634 4275 4708 4295
rect 4634 4223 4645 4275
rect 4697 4223 4708 4275
rect 4634 4185 4708 4223
rect 5150 4376 5224 4385
rect 5150 4320 5159 4376
rect 5215 4320 5224 4376
rect 5150 4295 5161 4320
rect 5213 4295 5224 4320
rect 5150 4275 5224 4295
rect 5150 4223 5161 4275
rect 5213 4223 5224 4275
rect 5150 4185 5224 4223
rect 5666 4376 5740 4385
rect 5666 4320 5675 4376
rect 5731 4320 5740 4376
rect 5666 4295 5677 4320
rect 5729 4295 5740 4320
rect 5666 4275 5740 4295
rect 5666 4223 5677 4275
rect 5729 4223 5740 4275
rect 5666 4185 5740 4223
rect 6293 4250 6373 4259
rect 6293 4194 6305 4250
rect 6361 4194 6373 4250
rect 6293 4183 6373 4194
rect 6505 4003 6585 4012
rect 6505 3947 6517 4003
rect 6573 3947 6585 4003
rect 6505 3936 6585 3947
rect 7630 3847 7676 4421
rect 8335 3799 8415 3808
rect 8335 3743 8347 3799
rect 8403 3743 8415 3799
rect 8335 3732 8415 3743
rect 10294 3672 10354 5675
rect 11071 4249 11200 4283
rect 11071 4193 11105 4249
rect 11161 4193 11200 4249
rect 11071 4161 11200 4193
rect 2891 3668 10354 3672
rect -2942 3616 10354 3668
rect 2916 3612 10354 3616
rect -2633 3561 -2553 3570
rect -2633 3505 -2621 3561
rect -2565 3505 -2553 3561
rect -2633 3494 -2553 3505
rect -2633 3283 -2553 3292
rect -2633 3227 -2621 3283
rect -2565 3227 -2553 3283
rect -2633 3216 -2553 3227
rect 7235 3274 7315 3283
rect 7235 3218 7247 3274
rect 7303 3218 7315 3274
rect 7235 3207 7315 3218
<< via2 >>
rect 2753 10903 2809 10959
rect 895 10412 951 10468
rect 3588 10661 3644 10690
rect 3588 10634 3590 10661
rect 3590 10634 3642 10661
rect 3642 10634 3644 10661
rect 4104 10537 4106 10562
rect 4106 10537 4158 10562
rect 4158 10537 4160 10562
rect 4104 10506 4160 10537
rect 4620 10661 4676 10690
rect 4620 10634 4622 10661
rect 4622 10634 4674 10661
rect 4674 10634 4676 10661
rect 9143 11083 9199 11139
rect 10022 11083 10078 11139
rect 3588 10119 3590 10142
rect 3590 10119 3642 10142
rect 3642 10119 3644 10142
rect 3588 10086 3644 10119
rect 4104 10243 4160 10271
rect 4104 10215 4106 10243
rect 4106 10215 4158 10243
rect 4158 10215 4160 10243
rect 4620 10119 4622 10141
rect 4622 10119 4674 10141
rect 4674 10119 4676 10141
rect 4620 10085 4676 10119
rect 3588 9825 3644 9854
rect 3588 9798 3590 9825
rect 3590 9798 3642 9825
rect 3642 9798 3644 9825
rect 4104 9701 4106 9724
rect 4106 9701 4158 9724
rect 4158 9701 4160 9724
rect 4104 9668 4160 9701
rect 4620 9825 4676 9854
rect 4620 9798 4622 9825
rect 4622 9798 4674 9825
rect 4674 9798 4676 9825
rect 3588 9283 3590 9306
rect 3590 9283 3642 9306
rect 3642 9283 3644 9306
rect 3588 9250 3644 9283
rect 4104 9407 4160 9435
rect 4104 9379 4106 9407
rect 4106 9379 4158 9407
rect 4158 9379 4160 9407
rect 4620 9283 4622 9306
rect 4622 9283 4674 9306
rect 4674 9283 4676 9306
rect 4620 9250 4676 9283
rect 3588 8985 3644 9014
rect 3588 8958 3590 8985
rect 3590 8958 3642 8985
rect 3642 8958 3644 8985
rect 4104 8861 4106 8883
rect 4106 8861 4158 8883
rect 4158 8861 4160 8883
rect 4104 8827 4160 8861
rect 4620 8985 4676 9014
rect 4620 8958 4622 8985
rect 4622 8958 4674 8985
rect 4674 8958 4676 8985
rect 3588 8439 3590 8462
rect 3590 8439 3642 8462
rect 3642 8439 3644 8462
rect 3588 8406 3644 8439
rect 4104 8563 4160 8592
rect 4104 8536 4106 8563
rect 4106 8536 4158 8563
rect 4158 8536 4160 8563
rect 4620 8439 4622 8462
rect 4622 8439 4674 8462
rect 4674 8439 4676 8462
rect 4620 8406 4676 8439
rect 2239 8371 2295 8374
rect 2239 8319 2241 8371
rect 2241 8319 2293 8371
rect 2293 8319 2295 8371
rect 2239 8318 2295 8319
rect -671 7912 -615 7941
rect -671 7885 -669 7912
rect -669 7885 -617 7912
rect -617 7885 -615 7912
rect -155 7912 -99 7941
rect -155 7885 -153 7912
rect -153 7885 -101 7912
rect -101 7885 -99 7912
rect 361 7912 417 7941
rect 361 7885 363 7912
rect 363 7885 415 7912
rect 415 7885 417 7912
rect 3209 7982 3265 7985
rect 3209 7930 3211 7982
rect 3211 7930 3263 7982
rect 3263 7930 3265 7982
rect 3209 7929 3265 7930
rect -1187 7494 -1131 7523
rect -1187 7467 -1185 7494
rect -1185 7467 -1133 7494
rect -1133 7467 -1131 7494
rect -671 7370 -669 7397
rect -669 7370 -617 7397
rect -617 7370 -615 7397
rect -671 7341 -615 7370
rect -155 7494 -99 7523
rect -155 7467 -153 7494
rect -153 7467 -101 7494
rect -101 7467 -99 7494
rect 361 7370 363 7397
rect 363 7370 415 7397
rect 415 7370 417 7397
rect 361 7341 417 7370
rect 877 7494 933 7523
rect 877 7467 879 7494
rect 879 7467 931 7494
rect 931 7467 933 7494
rect -1703 7076 -1647 7105
rect -1703 7049 -1701 7076
rect -1701 7049 -1649 7076
rect -1649 7049 -1647 7076
rect -1187 6952 -1185 6979
rect -1185 6952 -1133 6979
rect -1133 6952 -1131 6979
rect -1187 6923 -1131 6952
rect -671 7076 -615 7105
rect -671 7049 -669 7076
rect -669 7049 -617 7076
rect -617 7049 -615 7076
rect -155 6952 -153 6979
rect -153 6952 -101 6979
rect -101 6952 -99 6979
rect -155 6923 -99 6952
rect 361 7076 417 7105
rect 361 7049 363 7076
rect 363 7049 415 7076
rect 415 7049 417 7076
rect 877 6952 879 6979
rect 879 6952 931 6979
rect 931 6952 933 6979
rect 877 6923 933 6952
rect -1703 6534 -1701 6561
rect -1701 6534 -1649 6561
rect -1649 6534 -1647 6561
rect -1703 6505 -1647 6534
rect -1187 6658 -1131 6687
rect -1187 6631 -1185 6658
rect -1185 6631 -1133 6658
rect -1133 6631 -1131 6658
rect -671 6534 -669 6561
rect -669 6534 -617 6561
rect -617 6534 -615 6561
rect -671 6505 -615 6534
rect -155 6658 -99 6687
rect -155 6631 -153 6658
rect -153 6631 -101 6658
rect -101 6631 -99 6658
rect 361 6534 363 6561
rect 363 6534 415 6561
rect 415 6534 417 6561
rect 361 6505 417 6534
rect 877 6658 933 6687
rect 877 6631 879 6658
rect 879 6631 931 6658
rect 931 6631 933 6658
rect -1703 6240 -1647 6269
rect -1703 6213 -1701 6240
rect -1701 6213 -1649 6240
rect -1649 6213 -1647 6240
rect -1187 6116 -1185 6143
rect -1185 6116 -1133 6143
rect -1133 6116 -1131 6143
rect -1187 6087 -1131 6116
rect -671 6240 -615 6269
rect -671 6213 -669 6240
rect -669 6213 -617 6240
rect -617 6213 -615 6240
rect -155 6116 -153 6143
rect -153 6116 -101 6143
rect -101 6116 -99 6143
rect -155 6087 -99 6116
rect 361 6240 417 6269
rect 361 6213 363 6240
rect 363 6213 415 6240
rect 415 6213 417 6240
rect 877 6116 879 6143
rect 879 6116 931 6143
rect 931 6116 933 6143
rect 877 6087 933 6116
rect -1703 5698 -1701 5725
rect -1701 5698 -1649 5725
rect -1649 5698 -1647 5725
rect -1703 5669 -1647 5698
rect -1187 5822 -1131 5851
rect -1187 5795 -1185 5822
rect -1185 5795 -1133 5822
rect -1133 5795 -1131 5822
rect -671 5698 -669 5725
rect -669 5698 -617 5725
rect -617 5698 -615 5725
rect -671 5669 -615 5698
rect -155 5822 -99 5851
rect -155 5795 -153 5822
rect -153 5795 -101 5822
rect -101 5795 -99 5822
rect 361 5698 363 5725
rect 363 5698 415 5725
rect 415 5698 417 5725
rect 361 5669 417 5698
rect 877 5822 933 5851
rect 877 5795 879 5822
rect 879 5795 931 5822
rect 931 5795 933 5822
rect -1703 5404 -1647 5433
rect -1703 5377 -1701 5404
rect -1701 5377 -1649 5404
rect -1649 5377 -1647 5404
rect -1187 5280 -1185 5307
rect -1185 5280 -1133 5307
rect -1133 5280 -1131 5307
rect -1187 5251 -1131 5280
rect -671 5404 -615 5433
rect -671 5377 -669 5404
rect -669 5377 -617 5404
rect -617 5377 -615 5404
rect -155 5280 -153 5307
rect -153 5280 -101 5307
rect -101 5280 -99 5307
rect -155 5251 -99 5280
rect 361 5404 417 5433
rect 361 5377 363 5404
rect 363 5377 415 5404
rect 415 5377 417 5404
rect 877 5280 879 5307
rect 879 5280 931 5307
rect 931 5280 933 5307
rect 877 5251 933 5280
rect -1703 4862 -1701 4889
rect -1701 4862 -1649 4889
rect -1649 4862 -1647 4889
rect -1703 4833 -1647 4862
rect -1187 4986 -1131 5015
rect -1187 4959 -1185 4986
rect -1185 4959 -1133 4986
rect -1133 4959 -1131 4986
rect -671 4862 -669 4889
rect -669 4862 -617 4889
rect -617 4862 -615 4889
rect -671 4833 -615 4862
rect -155 4986 -99 5015
rect -155 4959 -153 4986
rect -153 4959 -101 4986
rect -101 4959 -99 4986
rect 361 4862 363 4889
rect 363 4862 415 4889
rect 415 4862 417 4889
rect 361 4833 417 4862
rect 877 4986 933 5015
rect 877 4959 879 4986
rect 879 4959 931 4986
rect 931 4959 933 4986
rect -1703 4568 -1647 4597
rect -1703 4541 -1701 4568
rect -1701 4541 -1649 4568
rect -1649 4541 -1647 4568
rect -1187 4444 -1185 4471
rect -1185 4444 -1133 4471
rect -1133 4444 -1131 4471
rect -1187 4415 -1131 4444
rect -671 4568 -615 4597
rect -671 4541 -669 4568
rect -669 4541 -617 4568
rect -617 4541 -615 4568
rect -155 4444 -153 4471
rect -153 4444 -101 4471
rect -101 4444 -99 4471
rect -155 4415 -99 4444
rect 361 4568 417 4597
rect 361 4541 363 4568
rect 363 4541 415 4568
rect 415 4541 417 4568
rect 4127 7273 4183 7302
rect 4127 7246 4129 7273
rect 4129 7246 4181 7273
rect 4181 7246 4183 7273
rect 4643 7273 4699 7302
rect 4643 7246 4645 7273
rect 4645 7246 4697 7273
rect 4697 7246 4699 7273
rect 5159 7273 5215 7302
rect 5159 7246 5161 7273
rect 5161 7246 5213 7273
rect 5213 7246 5215 7273
rect 5675 7273 5731 7302
rect 5675 7246 5677 7273
rect 5677 7246 5729 7273
rect 5729 7246 5731 7273
rect 4127 6855 4183 6884
rect 4127 6828 4129 6855
rect 4129 6828 4181 6855
rect 4181 6828 4183 6855
rect 4643 6731 4645 6758
rect 4645 6731 4697 6758
rect 4697 6731 4699 6758
rect 4643 6702 4699 6731
rect 5159 6855 5215 6884
rect 5159 6828 5161 6855
rect 5161 6828 5213 6855
rect 5213 6828 5215 6855
rect 5675 6731 5677 6758
rect 5677 6731 5729 6758
rect 5729 6731 5731 6758
rect 5675 6702 5731 6731
rect 4127 6313 4129 6340
rect 4129 6313 4181 6340
rect 4181 6313 4183 6340
rect 4127 6284 4183 6313
rect 4643 6437 4699 6466
rect 4643 6410 4645 6437
rect 4645 6410 4697 6437
rect 4697 6410 4699 6437
rect 5159 6313 5161 6340
rect 5161 6313 5213 6340
rect 5213 6313 5215 6340
rect 5159 6284 5215 6313
rect 5675 6437 5731 6466
rect 5675 6410 5677 6437
rect 5677 6410 5729 6437
rect 5729 6410 5731 6437
rect 4127 6019 4183 6048
rect 4127 5992 4129 6019
rect 4129 5992 4181 6019
rect 4181 5992 4183 6019
rect 4643 5895 4645 5922
rect 4645 5895 4697 5922
rect 4697 5895 4699 5922
rect 4643 5866 4699 5895
rect 5159 6019 5215 6048
rect 5159 5992 5161 6019
rect 5161 5992 5213 6019
rect 5213 5992 5215 6019
rect 5675 5895 5677 5922
rect 5677 5895 5729 5922
rect 5729 5895 5731 5922
rect 5675 5866 5731 5895
rect 4127 5477 4129 5504
rect 4129 5477 4181 5504
rect 4181 5477 4183 5504
rect 4127 5448 4183 5477
rect 4643 5601 4699 5630
rect 4643 5574 4645 5601
rect 4645 5574 4697 5601
rect 4697 5574 4699 5601
rect 5159 5477 5161 5504
rect 5161 5477 5213 5504
rect 5213 5477 5215 5504
rect 5159 5448 5215 5477
rect 5675 5601 5731 5630
rect 5675 5574 5677 5601
rect 5677 5574 5729 5601
rect 5729 5574 5731 5601
rect 4127 5183 4183 5212
rect 4127 5156 4129 5183
rect 4129 5156 4181 5183
rect 4181 5156 4183 5183
rect 4643 5059 4645 5086
rect 4645 5059 4697 5086
rect 4697 5059 4699 5086
rect 4643 5030 4699 5059
rect 5159 5183 5215 5212
rect 5159 5156 5161 5183
rect 5161 5156 5213 5183
rect 5213 5156 5215 5183
rect 5675 5059 5677 5086
rect 5677 5059 5729 5086
rect 5729 5059 5731 5086
rect 5675 5030 5731 5059
rect 4127 4641 4129 4668
rect 4129 4641 4181 4668
rect 4181 4641 4183 4668
rect 4127 4612 4183 4641
rect 4643 4765 4699 4794
rect 4643 4738 4645 4765
rect 4645 4738 4697 4765
rect 4697 4738 4699 4765
rect 5159 4641 5161 4668
rect 5161 4641 5213 4668
rect 5213 4641 5215 4668
rect 5159 4612 5215 4641
rect 5675 4765 5731 4794
rect 5675 4738 5677 4765
rect 5677 4738 5729 4765
rect 5729 4738 5731 4765
rect -1187 4150 -1131 4179
rect -1187 4123 -1185 4150
rect -1185 4123 -1133 4150
rect -1133 4123 -1131 4150
rect -671 4150 -615 4179
rect -671 4123 -669 4150
rect -669 4123 -617 4150
rect -617 4123 -615 4150
rect -155 4150 -99 4179
rect -155 4123 -153 4150
rect -153 4123 -101 4150
rect -101 4123 -99 4150
rect 1393 4050 1449 4053
rect 1393 3998 1395 4050
rect 1395 3998 1447 4050
rect 1447 3998 1449 4050
rect 1393 3997 1449 3998
rect 1507 4050 1563 4053
rect 1507 3998 1509 4050
rect 1509 3998 1561 4050
rect 1561 3998 1563 4050
rect 1507 3997 1563 3998
rect 4127 4347 4183 4376
rect 4127 4320 4129 4347
rect 4129 4320 4181 4347
rect 4181 4320 4183 4347
rect 4643 4347 4699 4376
rect 4643 4320 4645 4347
rect 4645 4320 4697 4347
rect 4697 4320 4699 4347
rect 5159 4347 5215 4376
rect 5159 4320 5161 4347
rect 5161 4320 5213 4347
rect 5213 4320 5215 4347
rect 5675 4347 5731 4376
rect 5675 4320 5677 4347
rect 5677 4320 5729 4347
rect 5729 4320 5731 4347
rect 6305 4247 6361 4250
rect 6305 4195 6307 4247
rect 6307 4195 6359 4247
rect 6359 4195 6361 4247
rect 6305 4194 6361 4195
rect 6517 4000 6573 4003
rect 6517 3948 6519 4000
rect 6519 3948 6571 4000
rect 6571 3948 6573 4000
rect 6517 3947 6573 3948
rect 8347 3796 8403 3799
rect 8347 3744 8349 3796
rect 8349 3744 8401 3796
rect 8401 3744 8403 3796
rect 8347 3743 8403 3744
rect 11105 4247 11161 4249
rect 11105 4195 11107 4247
rect 11107 4195 11159 4247
rect 11159 4195 11161 4247
rect 11105 4193 11161 4195
rect -2621 3558 -2565 3561
rect -2621 3506 -2619 3558
rect -2619 3506 -2567 3558
rect -2567 3506 -2565 3558
rect -2621 3505 -2565 3506
rect -2621 3280 -2565 3283
rect -2621 3228 -2619 3280
rect -2619 3228 -2567 3280
rect -2567 3228 -2565 3280
rect -2621 3227 -2565 3228
rect 7247 3271 7303 3274
rect 7247 3219 7249 3271
rect 7249 3219 7301 3271
rect 7301 3219 7303 3271
rect 7247 3218 7303 3219
<< metal3 >>
rect 915 11139 10087 11148
rect 915 11133 9143 11139
rect 886 11088 9143 11133
rect 886 10468 960 11088
rect 5850 11083 9143 11088
rect 9199 11083 10022 11139
rect 10078 11083 10087 11139
rect 5850 11074 10087 11083
rect 2744 10959 2818 10968
rect 2744 10903 2753 10959
rect 2809 10903 2818 10959
rect 2744 10699 2818 10903
rect 2610 10690 4685 10699
rect 2610 10634 3588 10690
rect 3644 10634 4620 10690
rect 4676 10634 4685 10690
rect 2610 10627 4685 10634
rect 886 10412 895 10468
rect 951 10412 960 10468
rect 886 10390 960 10412
rect 2744 10281 2818 10627
rect 5850 10567 5910 11074
rect 4095 10562 5910 10567
rect 4095 10506 4104 10562
rect 4160 10506 5910 10562
rect 4095 10495 5910 10506
rect 2610 10271 4169 10281
rect 2610 10215 4104 10271
rect 4160 10215 4169 10271
rect 2610 10209 4169 10215
rect 2744 9863 2818 10209
rect 5850 10148 5910 10495
rect 3579 10142 5910 10148
rect 3579 10086 3588 10142
rect 3644 10141 5910 10142
rect 3644 10086 4620 10141
rect 3579 10085 4620 10086
rect 4676 10085 5910 10141
rect 3579 10076 5910 10085
rect 2610 9854 4685 9863
rect 2610 9798 3588 9854
rect 3644 9798 4620 9854
rect 4676 9798 4685 9854
rect 2610 9791 4685 9798
rect 2744 9445 2818 9791
rect 5850 9730 5910 10076
rect 4095 9724 5910 9730
rect 4095 9668 4104 9724
rect 4160 9668 5910 9724
rect 4095 9658 5910 9668
rect 2610 9435 4169 9445
rect 2610 9379 4104 9435
rect 4160 9379 4169 9435
rect 2610 9373 4169 9379
rect 2744 9022 2818 9373
rect 5850 9312 5910 9658
rect 3579 9306 5910 9312
rect 3579 9250 3588 9306
rect 3644 9250 4620 9306
rect 4676 9250 5910 9306
rect 3579 9240 5910 9250
rect 2610 9014 4685 9022
rect 2610 8958 3588 9014
rect 3644 8958 4620 9014
rect 4676 8958 4685 9014
rect 2610 8950 4685 8958
rect 2744 8600 2818 8950
rect 5850 8889 5910 9240
rect 4095 8883 5910 8889
rect 4095 8827 4104 8883
rect 4160 8827 5910 8883
rect 4095 8817 5910 8827
rect 2610 8592 4169 8600
rect 2610 8536 4104 8592
rect 4160 8536 4169 8592
rect 2610 8528 4169 8536
rect 5850 8468 5910 8817
rect 3579 8462 5910 8468
rect 3579 8406 3588 8462
rect 3644 8406 4620 8462
rect 4676 8406 5910 8462
rect 2231 8374 2303 8405
rect 3579 8396 5910 8406
rect 2231 8318 2239 8374
rect 2295 8318 2303 8374
rect -2630 7950 -2556 8184
rect -2630 7941 426 7950
rect -2630 7885 -671 7941
rect -615 7885 -155 7941
rect -99 7885 361 7941
rect 417 7885 426 7941
rect -2630 7878 426 7885
rect -2630 7534 -2556 7878
rect -2630 7523 942 7534
rect -2630 7467 -1187 7523
rect -1131 7467 -155 7523
rect -99 7467 877 7523
rect 933 7467 942 7523
rect -2630 7462 942 7467
rect -2630 7116 -2556 7462
rect 2231 7402 2303 8318
rect -1712 7397 2303 7402
rect -1712 7341 -671 7397
rect -615 7341 361 7397
rect 417 7341 2303 7397
rect -1712 7330 2303 7341
rect -2630 7105 942 7116
rect -2630 7049 -1703 7105
rect -1647 7049 -671 7105
rect -615 7049 361 7105
rect 417 7049 942 7105
rect -2630 7044 942 7049
rect -2630 6698 -2556 7044
rect 2231 6984 2303 7330
rect -1712 6979 2303 6984
rect -1712 6923 -1187 6979
rect -1131 6923 -155 6979
rect -99 6923 877 6979
rect 933 6923 2303 6979
rect -1712 6912 2303 6923
rect -2630 6687 942 6698
rect -2630 6631 -1187 6687
rect -1131 6631 -155 6687
rect -99 6631 877 6687
rect 933 6631 942 6687
rect -2630 6626 942 6631
rect -2630 6280 -2556 6626
rect 2231 6566 2303 6912
rect -1712 6561 2303 6566
rect -1712 6505 -1703 6561
rect -1647 6505 -671 6561
rect -615 6505 361 6561
rect 417 6505 2303 6561
rect -1712 6494 2303 6505
rect -2630 6269 942 6280
rect -2630 6213 -1703 6269
rect -1647 6213 -671 6269
rect -615 6213 361 6269
rect 417 6213 942 6269
rect -2630 6208 942 6213
rect -2630 5862 -2556 6208
rect 2231 6148 2303 6494
rect -1712 6143 2303 6148
rect -1712 6087 -1187 6143
rect -1131 6087 -155 6143
rect -99 6087 877 6143
rect 933 6087 2303 6143
rect -1712 6076 2303 6087
rect -2630 5851 942 5862
rect -2630 5795 -1187 5851
rect -1131 5795 -155 5851
rect -99 5795 877 5851
rect 933 5795 942 5851
rect -2630 5790 942 5795
rect -2630 5444 -2556 5790
rect 2231 5730 2303 6076
rect -1712 5725 2303 5730
rect -1712 5669 -1703 5725
rect -1647 5669 -671 5725
rect -615 5669 361 5725
rect 417 5669 2303 5725
rect -1712 5658 2303 5669
rect -2630 5433 942 5444
rect -2630 5377 -1703 5433
rect -1647 5377 -671 5433
rect -615 5377 361 5433
rect 417 5377 942 5433
rect -2630 5372 942 5377
rect -2630 5026 -2556 5372
rect 2231 5312 2303 5658
rect -1712 5307 2303 5312
rect -1712 5251 -1187 5307
rect -1131 5251 -155 5307
rect -99 5251 877 5307
rect 933 5251 2303 5307
rect -1712 5240 2303 5251
rect -2630 5015 942 5026
rect -2630 4959 -1187 5015
rect -1131 4959 -155 5015
rect -99 4959 877 5015
rect 933 4959 942 5015
rect -2630 4954 942 4959
rect -2630 4608 -2556 4954
rect 2231 4894 2303 5240
rect -1712 4889 2303 4894
rect -1712 4833 -1703 4889
rect -1647 4833 -671 4889
rect -615 4833 361 4889
rect 417 4833 2303 4889
rect -1712 4822 2303 4833
rect -2630 4597 942 4608
rect -2630 4541 -1703 4597
rect -1647 4541 -671 4597
rect -615 4541 361 4597
rect 417 4541 942 4597
rect -2630 4536 942 4541
rect -2630 4190 -2556 4536
rect 2231 4476 2303 4822
rect -1712 4471 2303 4476
rect -1712 4415 -1187 4471
rect -1131 4415 -155 4471
rect -99 4415 2303 4471
rect -1712 4404 2303 4415
rect -2630 4179 942 4190
rect -2630 4123 -1187 4179
rect -1131 4123 -671 4179
rect -615 4123 -155 4179
rect -99 4123 942 4179
rect -2630 4118 942 4123
rect -2630 3561 -2556 4118
rect 2231 4064 2303 4404
rect 3200 7985 3274 8001
rect 3200 7929 3209 7985
rect 3265 7929 3274 7985
rect 3200 7311 3274 7929
rect 3200 7302 5740 7311
rect 3200 7246 4127 7302
rect 4183 7246 4643 7302
rect 4699 7246 5159 7302
rect 5215 7246 5675 7302
rect 5731 7246 5740 7302
rect 3200 7239 5740 7246
rect 3200 6895 3274 7239
rect 3200 6884 5740 6895
rect 3200 6828 4127 6884
rect 4183 6828 5159 6884
rect 5215 6828 5740 6884
rect 3200 6823 5740 6828
rect 3200 6477 3274 6823
rect 6508 6763 6580 7153
rect 4118 6758 6580 6763
rect 4118 6702 4643 6758
rect 4699 6702 5675 6758
rect 5731 6702 6580 6758
rect 4118 6691 6580 6702
rect 3200 6466 5740 6477
rect 3200 6410 4643 6466
rect 4699 6410 5675 6466
rect 5731 6410 5740 6466
rect 3200 6405 5740 6410
rect 3200 6059 3274 6405
rect 6508 6345 6580 6691
rect 4118 6340 6580 6345
rect 4118 6284 4127 6340
rect 4183 6284 5159 6340
rect 5215 6284 6580 6340
rect 4118 6273 6580 6284
rect 3200 6048 5740 6059
rect 3200 5992 4127 6048
rect 4183 5992 5159 6048
rect 5215 5992 5740 6048
rect 3200 5987 5740 5992
rect 3200 5641 3274 5987
rect 6508 5927 6580 6273
rect 4118 5922 6580 5927
rect 4118 5866 4643 5922
rect 4699 5866 5675 5922
rect 5731 5866 6580 5922
rect 4118 5855 6580 5866
rect 3200 5630 5740 5641
rect 3200 5574 4643 5630
rect 4699 5574 5675 5630
rect 5731 5574 5740 5630
rect 3200 5569 5740 5574
rect 3200 5223 3274 5569
rect 6508 5509 6580 5855
rect 4118 5504 6580 5509
rect 4118 5448 4127 5504
rect 4183 5448 5159 5504
rect 5215 5448 6580 5504
rect 4118 5437 6580 5448
rect 3200 5212 5740 5223
rect 3200 5156 4127 5212
rect 4183 5156 5159 5212
rect 5215 5156 5740 5212
rect 3200 5151 5740 5156
rect 3200 4805 3274 5151
rect 6508 5091 6580 5437
rect 4118 5086 6580 5091
rect 4118 5030 4643 5086
rect 4699 5030 5675 5086
rect 5731 5030 6580 5086
rect 4118 5019 6580 5030
rect 3200 4794 5740 4805
rect 3200 4738 4643 4794
rect 4699 4738 5675 4794
rect 5731 4738 5740 4794
rect 3200 4733 5740 4738
rect 3200 4387 3274 4733
rect 6508 4673 6580 5019
rect 4118 4668 6580 4673
rect 4118 4612 4127 4668
rect 4183 4612 5159 4668
rect 5215 4612 6580 4668
rect 4118 4601 6580 4612
rect 3200 4376 5740 4387
rect 3200 4320 4127 4376
rect 4183 4320 4643 4376
rect 4699 4320 5159 4376
rect 5215 4320 5675 4376
rect 5731 4320 5740 4376
rect 3200 4315 5740 4320
rect 3200 4314 3274 4315
rect 6508 4255 6580 4601
rect 4118 4250 6580 4255
rect 4118 4194 6305 4250
rect 6361 4194 6580 4250
rect 4118 4183 6580 4194
rect 1370 4053 2303 4064
rect 1370 3997 1393 4053
rect 1449 3997 1507 4053
rect 1563 3997 2303 4053
rect 1370 3984 2303 3997
rect 2231 3808 2303 3984
rect 6508 4003 6580 4183
rect 11071 4253 11200 4283
rect 11071 4189 11101 4253
rect 11165 4189 11200 4253
rect 11071 4161 11200 4189
rect 6508 3947 6517 4003
rect 6573 3947 6580 4003
rect 6508 3808 6580 3947
rect 2231 3799 12615 3808
rect 2231 3743 8347 3799
rect 8403 3743 12615 3799
rect 2231 3734 12615 3743
rect -2630 3505 -2621 3561
rect -2565 3505 -2556 3561
rect -2630 3465 -2556 3505
rect -2999 3283 -2200 3366
rect -2999 3227 -2621 3283
rect -2565 3227 -2200 3283
rect -2999 3184 -2200 3227
rect 6761 3274 7823 3338
rect 6761 3218 7247 3274
rect 7303 3218 7823 3274
rect 6761 3184 7823 3218
rect 10470 3184 11347 3190
rect -3733 -3896 11347 3184
<< via3 >>
rect 11101 4249 11165 4253
rect 11101 4193 11105 4249
rect 11105 4193 11161 4249
rect 11161 4193 11165 4249
rect 11101 4189 11165 4193
<< mimcap >>
rect -3693 3076 11307 3144
rect -3693 -3788 -3625 3076
rect 11239 -3788 11307 3076
rect -3693 -3856 11307 -3788
<< mimcapcontact >>
rect -3625 -3788 11239 3076
<< metal4 >>
rect 10200 4253 11273 4400
rect 10200 4189 11101 4253
rect 11165 4189 11273 4253
rect 10200 3104 11273 4189
rect -3653 3076 11273 3104
rect -3653 -3788 -3625 3076
rect 11239 2200 11273 3076
rect 11239 -3788 11267 2200
rect -3653 -3816 11267 -3788
use sky130_fd_pr__res_xhigh_po_1p41_THFN8M  sky130_fd_pr__res_xhigh_po_1p41_THFN8M_0
timestamp 1761058420
transform 1 0 10050 0 1 9377
box -297 -1672 297 1672
<< labels >>
flabel metal1 s 12197 11236 12197 11236 2 FreeSans 280 0 0 0 VDD
port 1 ne
flabel metal1 s 12012 8534 12012 8534 2 FreeSans 280 0 0 0 VOUT
port 5 ne
flabel metal2 s 12066 5701 12066 5701 2 FreeSans 280 0 0 0 IBIAS
port 2 ne
flabel metal2 s -4625 8653 -4625 8653 2 FreeSans 280 0 0 0 VN
port 3 ne
flabel metal2 s -4632 11141 -4632 11141 2 FreeSans 280 0 0 0 VP
port 4 ne
flabel metal2 s 11971 7303 11971 7303 2 FreeSans 280 0 0 0 EN
port 6 ne
flabel metal3 s 12161 3771 12161 3771 2 FreeSans 600 0 0 0 VSS
port 7 ne
<< properties >>
string FIXED_BBOX -3733 -3896 11347 3184
<< end >>
