** sch_path: /foss/designs/sky130_op_amp/runs/RUN_2025-10-21_16-29-21/parameters/dc_params/run_0/ac.sch
**.subckt ac
C1 Vout VSS {cl} m=1
Vdm net2 GND ac 1
Vcm net1 GND {vcm}
I0 VDD IBIAS {ib}
E2 VN net1 net2 GND -0.5
E1 VP net1 net2 GND 0.5
V0 VSS GND 0
V4 VDD GND {vdd}}
x1 VDD IBIAS VN VP Vout VDD VSS sky130_op_amp
**** begin user architecture code


.lib {PDK_ROOT}/{PDK}/libs.tech/combined/sky130.libs.spice {corner}

.include {DUT_path}

.temp {temperature}





.control
	* run ac simulation
	ac dec 20 1k 100e6

	* measure parameters
	let vout_mag = abs(v(Vout))
	let vout_phase_margin = phase(v(Vout)) * 180/pi + 180
	meas ac A0 find vout_mag at=1k
	meas ac UGF when vout_mag=1 fall=1
	meas ac PM find vout_phase_margin when vout_mag=1

	echo $&A0 $&ugf $&PM > {simpath}/{filename}_{N}.data
	quit
.endc



**** end user architecture code
**.ends
.GLOBAL GND
.end
