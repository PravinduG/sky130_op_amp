** sch_path: /foss/designs/sky130_op_amp/runs/RUN_2025-10-22_16-40-42/parameters/dc_params/run_44/sky130_op_amp_tb.sch
**.subckt sky130_op_amp_tb
C1 Vout VSS 2.5e-11 m=1
Vdm net2 GND ac 1
Vcm net1 GND 0.9
I0 VDD IBIAS 4.9999999999999996e-06
E2 VN net1 net2 GND -0.5
E1 VP net1 net2 GND 0.5
V0 VSS GND 0
V4 VDD GND 1.9
x1 VDD IBIAS VN VP Vout VDD VSS sky130_op_amp
**** begin user architecture code


.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice sf

.include /foss/designs/sky130_op_amp/netlist/rcx/sky130_op_amp.spice

.temp 50

.option SEED=12345

* Flag unsafe operating conditions (exceeds models' specified limits)
.option warn=1




.control
	* run ac simulation
	ac dec 20 1k 100e6

	* measure parameters
	let vout_mag = dB(abs(v(Vout)))
	let vout_phase_margin = phase(v(Vout)) * 180/pi + 180
	meas ac A0 find vout_mag at=1k
	meas ac UGF when vout_mag=1 fall=1
	meas ac PM find vout_phase_margin when vout_mag=1

	echo $&A0 $&ugf $&PM > /foss/designs/sky130_op_amp/runs/RUN_2025-10-22_16-40-42/parameters/dc_params/run_44/sky130_op_amp_tb_44.data
.endc



**** end user architecture code
**.ends
.GLOBAL GND
.end
