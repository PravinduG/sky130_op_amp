* NGSPICE file created from sky130_op_amp.ext - technology: sky130A

.subckt sky130_op_amp VDD IBIAS VN VP VOUT EN VSS
X0 a_8862_4192.t27 EN.t0 VSS.t311 VSS.t215 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1 VDD.t97 VDD.t96 VDD.t97 VDD.t44 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X2 VDD.t95 VDD.t93 VDD.t94 VDD.t47 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X3 a_3868_4185.t39 IBIAS.t10 a_3329_8823.t39 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X4 a_n1962_4406.t59 IBIAS.t11 VOUT.t21 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X5 a_n1962_4406.t58 IBIAS.t12 VOUT.t53 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X6 VSS.t211 VSS.t209 VSS.t210 VSS.t30 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X7 a_3329_8823.t38 IBIAS.t13 a_3868_4185.t38 VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X8 VSS.t208 VSS.t207 VSS.t208 VSS.t64 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X9 VDD.t92 VDD.t91 VDD.t92 VDD.t71 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X10 a_3868_4185.t37 IBIAS.t14 a_3329_8823.t8 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X11 a_n735_8972.t23 VP.t0 a_3329_8823.t56 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X12 VSS.t310 EN.t1 a_n1962_4406.t123 VSS.t77 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X13 a_3868_4185.t36 IBIAS.t15 a_3329_8823.t17 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X14 a_3329_8823.t66 VN.t0 a_n935_8875.t15 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X15 VDD.t19 a_n735_8972.t27 VOUT.t67 VDD.t15 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X16 a_n1962_4406.t122 EN.t2 VSS.t309 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X17 a_3329_8823.t65 VN.t1 a_n935_8875.t14 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X18 VDD.t36 a_n735_8972.t28 VOUT.t77 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X19 VSS.t206 VSS.t205 a_3329_8823.t55 VSS.t64 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X20 a_n1962_4406.t57 IBIAS.t16 VOUT.t45 VSS.t212 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X21 a_n1962_4406.t56 IBIAS.t17 VOUT.t2 VSS.t212 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X22 VSS.t308 EN.t3 a_n1962_4406.t121 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X23 a_3329_8823.t43 VN.t2 a_n935_8875.t13 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X24 VDD.t90 VDD.t89 VDD.t90 VDD.t71 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X25 a_n1962_4406.t79 VSS.t203 VSS.t204 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X26 a_n1962_4406.t120 EN.t4 VSS.t307 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X27 VOUT.t38 IBIAS.t18 a_n1962_4406.t55 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X28 VSS.t202 VSS.t201 a_n1962_4406.t78 VSS.t56 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X29 VDD.t88 VDD.t87 VDD.t88 VDD.t44 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X30 a_n935_8875.t12 VN.t3 a_3329_8823.t62 VSS.t84 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X31 VOUT.t46 IBIAS.t19 a_n1962_4406.t54 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X32 VDD.t86 VDD.t84 VDD.t85 VDD.t47 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X33 a_3329_8823.t63 VP.t1 a_n735_8972.t22 VSS.t89 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X34 VSS.t306 EN.t5 a_n1962_4406.t119 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X35 VDD.t17 a_n735_8972.t29 VOUT.t65 VDD.t15 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X36 VDD.t16 a_n735_8972.t30 VOUT.t64 VDD.t15 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X37 VSS.t198 VSS.t197 VSS.t198 VSS.t56 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X38 a_n1962_4406.t53 IBIAS.t20 VOUT.t42 VSS.t45 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X39 VOUT.t35 IBIAS.t21 a_n1962_4406.t52 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X40 VSS.t200 VSS.t199 a_3868_4185.t55 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X41 VSS.t196 VSS.t195 a_3868_4185.t54 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X42 a_n1962_4406.t77 VSS.t193 VSS.t194 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X43 a_3329_8823.t42 VN.t4 a_n935_8875.t11 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X44 a_n1962_4406.t118 EN.t6 VSS.t305 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X45 a_n1962_4406.t117 EN.t7 VSS.t304 VSS.t212 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X46 VSS.t192 VSS.t191 VSS.t192 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X47 a_n735_8972.t21 VP.t2 a_3329_8823.t73 VSS.t313 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X48 a_n1962_4406.t51 IBIAS.t22 VOUT.t9 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X49 a_n1962_4406.t116 EN.t8 VSS.t303 VSS.t212 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X50 a_3329_8823.t35 IBIAS.t23 a_3868_4185.t35 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X51 IBIAS.t7 IBIAS.t6 a_8862_4192.t0 VSS.t214 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X52 VSS.t302 EN.t9 a_8862_4192.t26 VSS.t214 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X53 a_n935_8875.t33 a_n935_8875.t32 VDD.t110 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X54 a_n1962_4406.t50 IBIAS.t24 VOUT.t3 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X55 VSS.t190 VSS.t188 VSS.t189 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X56 VOUT.t0 IBIAS.t25 a_n1962_4406.t49 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X57 VOUT.t6 IBIAS.t26 a_n1962_4406.t48 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X58 a_3868_4185.t53 VSS.t186 VSS.t187 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X59 a_8862_4192.t25 EN.t10 VSS.t301 VSS.t219 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X60 VSS.t185 VSS.t183 VSS.t184 VSS.t30 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X61 VDD.t7 a_n735_8972.t31 VOUT.t62 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X62 a_n735_8972.t7 a_9909_7861.t0 VSS.t218 sky130_fd_pr__res_xhigh_po_1p41 l=11
X63 a_3868_4185.t34 IBIAS.t27 a_3329_8823.t4 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X64 a_8862_4192.t3 IBIAS.t4 IBIAS.t5 VSS.t219 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X65 VSS.t300 EN.t11 a_n1962_4406.t115 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X66 a_n1962_4406.t114 EN.t12 VSS.t299 VSS.t45 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X67 VSS.t182 VSS.t181 VSS.t182 VSS.t45 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X68 a_n735_8972.t24 a_n935_8875.t34 VDD.t103 VDD.t30 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X69 VSS.t180 VSS.t179 a_3329_8823.t54 VSS.t64 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X70 a_3329_8823.t2 IBIAS.t28 a_3868_4185.t33 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X71 VSS.t178 VSS.t177 VSS.t178 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X72 VSS.t293 EN.t13 a_3868_4185.t79 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X73 a_n935_8875.t10 VN.t5 a_3329_8823.t64 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X74 VSS.t298 EN.t14 a_n1962_4406.t113 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X75 VSS.t176 VSS.t175 a_n1962_4406.t76 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X76 a_3329_8823.t71 VN.t6 a_n935_8875.t9 VSS.t89 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X77 VDD.t83 VDD.t82 VDD.t83 VDD.t71 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X78 a_3868_4185.t78 EN.t15 VSS.t297 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X79 a_3868_4185.t77 EN.t16 VSS.t296 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X80 VDD.t33 a_n735_8972.t32 VOUT.t75 VDD.t15 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X81 VSS.t295 EN.t17 a_8862_4192.t24 VSS.t214 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X82 a_3329_8823.t28 IBIAS.t29 a_3868_4185.t32 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X83 a_3329_8823.t77 VP.t3 a_n735_8972.t20 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X84 VDD.t105 a_n735_8972.t33 VOUT.t86 VDD.t15 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X85 a_3868_4185.t31 IBIAS.t30 a_3329_8823.t11 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X86 a_n1962_4406.t112 EN.t18 VSS.t294 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X87 a_8862_4192.t23 EN.t19 VSS.t292 VSS.t219 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X88 VSS.t174 VSS.t172 VSS.t173 VSS.t30 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X89 a_3329_8823.t12 IBIAS.t31 a_3868_4185.t30 VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X90 a_3868_4185.t52 VSS.t170 VSS.t171 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X91 VOUT.t49 IBIAS.t32 a_n1962_4406.t47 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X92 VOUT.t28 IBIAS.t33 a_n1962_4406.t46 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X93 a_n1962_4406.t45 IBIAS.t34 VOUT.t57 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X94 a_3868_4185.t76 EN.t20 VSS.t291 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X95 a_3329_8823.t61 VP.t4 a_n735_8972.t19 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X96 VOUT.t69 a_n735_8972.t34 VDD.t23 VDD.t13 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X97 VSS.t130 VSS.t129 VSS.t130 VSS.t77 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X98 a_3868_4185.t75 EN.t21 VSS.t290 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X99 VSS.t289 EN.t22 a_3868_4185.t74 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X100 VOUT.t54 IBIAS.t35 a_n1962_4406.t44 VSS.t77 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X101 a_3868_4185.t29 IBIAS.t36 a_3329_8823.t18 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X102 VSS.t169 VSS.t168 VSS.t169 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X103 a_n1962_4406.t43 IBIAS.t37 VOUT.t52 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X104 VOUT.t25 IBIAS.t38 a_n1962_4406.t42 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X105 VSS.t167 VSS.t166 VSS.t167 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X106 VOUT.t26 IBIAS.t39 a_n1962_4406.t41 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X107 VSS.t165 VSS.t164 a_n1962_4406.t75 VSS.t56 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X108 VSS.t288 EN.t23 a_n1962_4406.t111 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X109 a_n935_8875.t8 VN.t7 a_3329_8823.t46 VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X110 VDD.t81 VDD.t80 VDD.t81 VDD.t71 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X111 VSS.t287 EN.t24 a_n1962_4406.t110 VSS.t77 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X112 VSS.t286 EN.t25 a_n1962_4406.t109 VSS.t77 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X113 VDD.t106 a_n935_8875.t35 a_n735_8972.t25 VDD.t11 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X114 a_n1962_4406.t40 IBIAS.t40 VOUT.t58 VSS.t45 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X115 VSS.t163 VSS.t161 VSS.t163 VSS.t162 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X116 VDD.t25 a_n735_8972.t35 VOUT.t71 VDD.t15 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X117 VSS.t160 VSS.t158 VSS.t159 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X118 a_n1962_4406.t108 EN.t26 VSS.t285 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X119 a_3329_8823.t27 IBIAS.t41 a_3868_4185.t28 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X120 a_n935_8875.t31 a_n935_8875.t30 VDD.t37 VDD.t30 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X121 a_n1962_4406.t39 IBIAS.t42 VOUT.t13 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X122 VOUT.t16 IBIAS.t43 a_n1962_4406.t38 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X123 a_n1962_4406.t37 IBIAS.t44 VOUT.t22 VSS.t212 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X124 a_n1962_4406.t107 EN.t27 VSS.t284 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X125 a_3329_8823.t0 IBIAS.t45 a_3868_4185.t27 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X126 a_n735_8972.t18 VP.t5 a_3329_8823.t47 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X127 VSS.t157 VSS.t155 a_n735_8972.t4 VSS.t156 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X128 VOUT.t73 a_n735_8972.t36 VDD.t27 VDD.t13 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X129 a_n1962_4406.t36 IBIAS.t46 VOUT.t39 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X130 a_n1962_4406.t106 EN.t28 VSS.t280 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X131 VSS.t281 EN.t29 a_n1962_4406.t105 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X132 VSS.t283 EN.t30 a_n1962_4406.t104 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X133 VSS.t282 EN.t31 a_8862_4192.t22 VSS.t214 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X134 a_3329_8823.t53 VSS.t153 VSS.t154 VSS.t61 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X135 VOUT.t14 IBIAS.t47 a_n1962_4406.t35 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X136 VSS.t152 VSS.t151 a_n1962_4406.t74 VSS.t56 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X137 VOUT.t17 IBIAS.t48 a_n1962_4406.t34 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X138 VSS.t150 VSS.t149 VSS.t150 VSS.t56 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X139 VSS.t279 EN.t32 a_n1962_4406.t103 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X140 a_n1962_4406.t33 IBIAS.t49 VOUT.t50 VSS.t212 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X141 a_3868_4185.t73 EN.t33 VSS.t278 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X142 VSS.t274 EN.t34 a_3868_4185.t72 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X143 VSS.t277 EN.t35 a_3868_4185.t71 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X144 a_n935_8875.t29 a_n935_8875.t28 VDD.t29 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X145 VDD.t79 VDD.t78 VDD.t79 VDD.t71 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X146 a_n1962_4406.t32 IBIAS.t50 VOUT.t29 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X147 a_8862_4192.t21 EN.t36 VSS.t276 VSS.t219 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X148 a_3868_4185.t70 EN.t37 VSS.t275 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X149 VSS.t148 VSS.t147 a_3868_4185.t51 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X150 VDD.t22 a_n935_8875.t26 a_n935_8875.t27 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X151 VOUT.t23 IBIAS.t51 a_n1962_4406.t31 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X152 VSS.t273 EN.t38 a_3868_4185.t69 VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X153 a_3868_4185.t50 VSS.t145 VSS.t146 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X154 VSS.t144 VSS.t142 VSS.t143 VSS.t30 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X155 a_3868_4185.t49 VSS.t140 VSS.t141 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X156 VSS.t272 EN.t39 a_3868_4185.t68 VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X157 VSS.t271 EN.t40 a_n1962_4406.t102 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X158 a_3868_4185.t26 IBIAS.t52 a_3329_8823.t14 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X159 a_3868_4185.t25 IBIAS.t53 a_3329_8823.t24 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X160 a_3329_8823.t67 VN.t8 a_n935_8875.t7 VSS.t217 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X161 a_3868_4185.t24 IBIAS.t54 a_3329_8823.t34 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X162 VDD.t77 VDD.t76 VDD.t77 VDD.t71 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X163 a_n1962_4406.t73 VSS.t138 VSS.t139 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X164 a_n1962_4406.t72 VSS.t136 VSS.t137 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X165 IBIAS.t3 IBIAS.t2 a_8862_4192.t2 VSS.t216 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X166 VSS.t270 EN.t41 a_8862_4192.t20 VSS.t216 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X167 a_3868_4185.t23 IBIAS.t55 a_3329_8823.t5 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X168 a_3329_8823.t9 IBIAS.t56 a_3868_4185.t22 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X169 a_n1962_4406.t101 EN.t42 VSS.t269 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X170 a_n1962_4406.t100 EN.t43 VSS.t268 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X171 a_3329_8823.t13 IBIAS.t57 a_3868_4185.t21 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X172 VDD.t75 VDD.t73 VDD.t74 VDD.t40 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X173 VSS.t267 EN.t44 a_8862_4192.t19 VSS.t214 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X174 a_8862_4192.t18 EN.t45 VSS.t266 VSS.t215 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X175 VDD.t101 a_n735_8972.t37 VOUT.t83 VDD.t15 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X176 a_n1962_4406.t30 IBIAS.t58 VOUT.t55 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X177 a_8862_4192.t1 IBIAS.t0 IBIAS.t1 VSS.t215 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X178 a_3329_8823.t1 IBIAS.t59 a_3868_4185.t20 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X179 VDD.t109 a_n935_8875.t36 a_n735_8972.t26 VDD.t11 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X180 a_8862_4192.t17 EN.t46 VSS.t265 VSS.t219 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X181 VSS.t135 VSS.t133 VSS.t134 VSS.t30 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X182 VOUT.t81 a_n735_8972.t38 VDD.t99 VDD.t13 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X183 VSS.t128 VSS.t127 a_3868_4185.t48 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X184 a_3868_4185.t47 VSS.t131 VSS.t132 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X185 a_n935_8875.t25 a_n935_8875.t24 VDD.t31 VDD.t30 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X186 a_3868_4185.t19 IBIAS.t60 a_3329_8823.t25 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X187 a_3329_8823.t52 VSS.t125 VSS.t126 VSS.t61 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X188 VSS.t248 EN.t47 a_8862_4192.t16 VSS.t216 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X189 a_3329_8823.t6 IBIAS.t61 a_3868_4185.t18 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X190 VDD.t72 VDD.t70 VDD.t72 VDD.t71 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X191 a_3868_4185.t67 EN.t48 VSS.t264 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X192 VOUT.t63 a_n735_8972.t39 VDD.t14 VDD.t13 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X193 VOUT.t68 a_n735_8972.t40 VDD.t20 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X194 a_n1962_4406.t99 EN.t49 VSS.t263 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X195 a_8862_4192.t15 EN.t50 VSS.t262 VSS.t215 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X196 VSS.t124 VSS.t123 a_3329_8823.t51 VSS.t64 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X197 a_n1962_4406.t98 EN.t51 VSS.t261 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X198 VDD.t69 VDD.t67 VDD.t68 VDD.t40 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X199 a_3329_8823.t58 VP.t6 a_n735_8972.t17 VSS.t89 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X200 VSS.t122 VSS.t121 a_n1962_4406.t71 VSS.t56 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X201 a_3329_8823.t79 VN.t9 a_n935_8875.t6 VSS.t89 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X202 VOUT.t40 IBIAS.t62 a_n1962_4406.t29 VSS.t77 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X203 a_n935_8875.t5 VN.t10 a_3329_8823.t70 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X204 VDD.t66 VDD.t64 VDD.t65 VDD.t40 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X205 a_n735_8972.t5 a_n935_8875.t37 VDD.t28 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X206 VOUT.t66 a_n735_8972.t41 VDD.t18 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X207 VSS.t120 VSS.t119 VSS.t120 VSS.t45 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X208 a_n1962_4406.t97 EN.t52 VSS.t260 VSS.t45 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X209 a_n1962_4406.t28 IBIAS.t63 VOUT.t15 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X210 VSS.t118 VSS.t117 VSS.t118 VSS.t77 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X211 VDD.t4 a_n935_8875.t38 a_n735_8972.t0 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X212 a_n735_8972.t16 VP.t7 a_3329_8823.t74 VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X213 a_3329_8823.t75 VP.t8 a_n735_8972.t15 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X214 a_n1962_4406.t96 EN.t53 VSS.t259 VSS.t212 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X215 VDD.t63 VDD.t61 VDD.t62 VDD.t40 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X216 VSS.t116 VSS.t115 a_n1962_4406.t70 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X217 a_n1962_4406.t27 IBIAS.t64 VOUT.t18 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X218 VSS.t258 EN.t54 a_n1962_4406.t95 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X219 VOUT.t10 IBIAS.t65 a_n1962_4406.t26 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X220 a_n735_8972.t14 VP.t9 a_3329_8823.t78 VSS.t84 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X221 a_3329_8823.t59 VP.t10 a_n735_8972.t13 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X222 a_n735_8972.t12 VP.t11 a_3329_8823.t69 VSS.t84 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X223 a_n1962_4406.t69 VSS.t113 VSS.t114 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X224 VSS.t257 EN.t55 a_n1962_4406.t94 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X225 a_n1962_4406.t68 VSS.t111 VSS.t112 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X226 VOUT.t51 IBIAS.t66 a_n1962_4406.t25 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X227 VOUT.t30 IBIAS.t67 a_n1962_4406.t24 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X228 VOUT.t24 IBIAS.t68 a_n1962_4406.t23 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X229 VSS.t256 EN.t56 a_8862_4192.t14 VSS.t214 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X230 a_8862_4192.t13 EN.t57 VSS.t255 VSS.t219 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X231 VDD.t21 a_n935_8875.t22 a_n935_8875.t23 VDD.t11 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X232 a_3329_8823.t50 VSS.t109 VSS.t110 VSS.t61 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X233 VOUT.t56 IBIAS.t69 a_n1962_4406.t22 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X234 a_n1962_4406.t21 IBIAS.t70 VOUT.t20 VSS.t45 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X235 a_3329_8823.t16 IBIAS.t71 a_3868_4185.t17 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X236 VSS.t108 VSS.t107 a_3868_4185.t46 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X237 VOUT.t79 a_n735_8972.t42 VDD.t38 VDD.t13 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X238 VOUT.t34 IBIAS.t72 a_n1962_4406.t20 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X239 a_n1962_4406.t19 IBIAS.t73 VOUT.t11 VSS.t45 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X240 VSS.t106 VSS.t105 a_3868_4185.t45 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X241 VSS.t104 VSS.t101 VSS.t103 VSS.t102 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X242 a_n1962_4406.t18 IBIAS.t74 VOUT.t31 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X243 VSS.t100 VSS.t99 VSS.t100 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X244 VSS.t254 EN.t58 a_8862_4192.t12 VSS.t216 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X245 VOUT.t8 IBIAS.t75 a_n1962_4406.t17 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X246 a_n1962_4406.t16 IBIAS.t76 VOUT.t32 VSS.t212 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X247 a_n1962_4406.t15 IBIAS.t77 VOUT.t4 VSS.t212 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X248 a_3868_4185.t16 IBIAS.t78 a_3329_8823.t21 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X249 VSS.t98 VSS.t97 IBIAS.t9 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X250 a_n1962_4406.t93 EN.t59 VSS.t253 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X251 VOUT.t19 IBIAS.t79 a_n1962_4406.t14 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X252 a_n1962_4406.t92 EN.t60 VSS.t252 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X253 a_3868_4185.t15 IBIAS.t80 a_3329_8823.t36 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X254 VSS.t251 EN.t61 a_8862_4192.t11 VSS.t214 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X255 VDD.t60 VDD.t58 VDD.t59 VDD.t47 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X256 a_n735_8972.t11 VP.t12 a_3329_8823.t40 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X257 VSS.t250 EN.t62 a_n1962_4406.t91 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X258 VSS.t96 VSS.t95 VSS.t96 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X259 a_8862_4192.t10 EN.t63 VSS.t249 VSS.t215 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X260 a_3868_4185.t14 IBIAS.t81 a_3329_8823.t32 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X261 VSS.t247 EN.t64 a_n1962_4406.t90 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X262 a_3329_8823.t23 IBIAS.t82 a_3868_4185.t13 VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X263 a_8862_4192.t9 EN.t65 VSS.t246 VSS.t219 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X264 VSS.t245 EN.t66 a_3868_4185.t66 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X265 a_n735_8972.t1 a_n935_8875.t39 VDD.t9 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X266 VDD.t35 a_n735_8972.t43 VOUT.t76 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X267 a_n1962_4406.t13 IBIAS.t83 VOUT.t43 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X268 a_3329_8823.t45 VN.t11 a_n935_8875.t4 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X269 VOUT.t88 a_n735_8972.t44 VDD.t108 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X270 VSS.t244 EN.t67 a_n1962_4406.t89 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X271 a_3868_4185.t12 IBIAS.t84 a_3329_8823.t10 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X272 VSS.t94 VSS.t93 a_3868_4185.t44 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X273 a_3868_4185.t43 VSS.t91 VSS.t92 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X274 a_3329_8823.t7 IBIAS.t85 a_3868_4185.t11 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X275 VDD.t10 a_n935_8875.t40 a_n735_8972.t2 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X276 VSS.t90 VSS.t88 a_n935_8875.t17 VSS.t89 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X277 a_n935_8875.t3 VN.t12 a_3329_8823.t57 VSS.t84 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X278 VDD.t57 VDD.t55 VDD.t56 VDD.t40 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X279 VSS.t243 EN.t68 a_n1962_4406.t88 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X280 a_3868_4185.t10 IBIAS.t86 a_3329_8823.t3 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X281 VSS.t87 VSS.t86 VSS.t87 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X282 VSS.t242 EN.t69 a_8862_4192.t8 VSS.t216 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X283 a_3329_8823.t29 IBIAS.t87 a_3868_4185.t9 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X284 VOUT.t74 a_n735_8972.t45 VDD.t32 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X285 a_3868_4185.t65 EN.t70 VSS.t241 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X286 VDD.t102 a_n735_8972.t46 VOUT.t84 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X287 a_8862_4192.t7 EN.t71 VSS.t240 VSS.t215 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X288 VSS.t239 EN.t72 a_3868_4185.t64 VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X289 VDD.t12 a_n935_8875.t20 a_n935_8875.t21 VDD.t11 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X290 a_n935_8875.t2 VN.t13 a_3329_8823.t68 VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X291 VDD.t54 VDD.t53 VDD.t54 VDD.t44 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X292 a_n935_8875.t16 VSS.t83 VSS.t85 VSS.t84 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X293 VSS.t82 VSS.t81 VSS.t82 VSS.t56 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X294 VOUT.t85 a_n735_8972.t47 VDD.t104 VDD.t13 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X295 VSS.t80 VSS.t79 a_n1962_4406.t67 VSS.t56 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X296 a_3868_4185.t8 IBIAS.t88 a_3329_8823.t26 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X297 VSS.t78 VSS.t76 VSS.t78 VSS.t77 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X298 VDD.t107 a_n735_8972.t48 VOUT.t87 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X299 a_n1962_4406.t66 VSS.t74 VSS.t75 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X300 VSS.t73 VSS.t71 VSS.t72 VSS.t61 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X301 VDD.t24 a_n735_8972.t49 VOUT.t70 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X302 VSS.t238 EN.t73 a_n1962_4406.t87 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X303 VSS.t70 VSS.t68 VSS.t69 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X304 VOUT.t72 a_n735_8972.t50 VDD.t26 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X305 VOUT.t41 IBIAS.t89 a_n1962_4406.t12 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X306 a_n1962_4406.t65 VSS.t66 VSS.t67 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X307 a_n1962_4406.t86 EN.t74 VSS.t237 VSS.t212 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X308 VSS.t65 VSS.t63 a_3329_8823.t49 VSS.t64 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X309 a_3329_8823.t48 VSS.t60 VSS.t62 VSS.t61 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X310 a_n1962_4406.t11 IBIAS.t90 VOUT.t47 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X311 VSS.t59 VSS.t58 a_n1962_4406.t64 VSS.t56 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X312 VDD.t1 a_n935_8875.t18 a_n935_8875.t19 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X313 a_n735_8972.t10 VP.t13 a_3329_8823.t41 VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X314 a_n935_8875.t1 VN.t14 a_3329_8823.t72 VSS.t312 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X315 VDD.t52 VDD.t50 VDD.t51 VDD.t40 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X316 VOUT.t44 IBIAS.t91 a_n1962_4406.t10 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X317 VSS.t57 VSS.t55 a_n1962_4406.t63 VSS.t56 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X318 a_3329_8823.t30 IBIAS.t92 a_3868_4185.t7 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X319 VDD.t49 VDD.t46 VDD.t48 VDD.t47 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X320 VOUT.t82 a_n735_8972.t51 VDD.t100 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X321 VOUT.t36 IBIAS.t93 a_n1962_4406.t9 VSS.t77 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X322 VOUT.t37 IBIAS.t94 a_n1962_4406.t8 VSS.t77 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X323 a_3329_8823.t22 IBIAS.t95 a_3868_4185.t6 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X324 a_3329_8823.t60 VP.t14 a_n735_8972.t9 VSS.t213 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X325 a_n1962_4406.t85 EN.t75 VSS.t236 VSS.t45 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X326 a_9909_7861.t1 VOUT.t78 sky130_fd_pr__cap_mim_m3_1 l=35 w=75
X327 a_3868_4185.t42 VSS.t53 VSS.t54 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X328 VOUT.t80 a_n735_8972.t52 VDD.t98 VDD.t13 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X329 a_n1962_4406.t7 IBIAS.t96 VOUT.t12 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X330 a_n1962_4406.t6 IBIAS.t97 VOUT.t5 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X331 a_3868_4185.t63 EN.t76 VSS.t235 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X332 VSS.t234 EN.t77 a_3868_4185.t62 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X333 VSS.t233 EN.t78 a_3868_4185.t61 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X334 a_3868_4185.t41 VSS.t50 VSS.t52 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X335 a_n735_8972.t6 a_n935_8875.t41 VDD.t34 VDD.t30 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X336 a_n735_8972.t3 VSS.t47 VSS.t49 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X337 a_n1962_4406.t84 EN.t79 VSS.t223 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X338 VSS.t232 EN.t80 a_n1962_4406.t83 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X339 VOUT.t1 IBIAS.t98 a_n1962_4406.t5 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X340 VSS.t46 VSS.t44 VSS.t46 VSS.t45 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X341 VSS.t43 VSS.t42 VSS.t43 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X342 a_3868_4185.t60 EN.t81 VSS.t231 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X343 a_3329_8823.t76 VP.t15 a_n735_8972.t8 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X344 a_n1962_4406.t62 VSS.t40 VSS.t41 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X345 VSS.t228 EN.t82 a_n1962_4406.t82 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X346 VOUT.t7 IBIAS.t99 a_n1962_4406.t4 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X347 a_n1962_4406.t61 VSS.t37 VSS.t39 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X348 VSS.t230 EN.t83 a_n1962_4406.t81 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X349 VSS.t229 EN.t84 a_3868_4185.t59 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X350 VSS.t227 EN.t85 a_8862_4192.t6 VSS.t216 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X351 VSS.t226 EN.t86 a_3868_4185.t58 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X352 VSS.t36 VSS.t35 VSS.t36 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X353 a_3868_4185.t5 IBIAS.t100 a_3329_8823.t15 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X354 a_3868_4185.t4 IBIAS.t101 a_3329_8823.t37 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X355 a_n1962_4406.t3 IBIAS.t102 VOUT.t48 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X356 a_8862_4192.t5 EN.t87 VSS.t225 VSS.t215 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X357 VOUT.t60 a_n735_8972.t53 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X358 VDD.t6 a_n735_8972.t54 VOUT.t61 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X359 a_n1962_4406.t80 EN.t88 VSS.t224 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X360 a_3329_8823.t33 IBIAS.t103 a_3868_4185.t3 VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X361 IBIAS.t8 VSS.t33 VSS.t34 VSS.t30 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X362 VSS.t32 VSS.t29 VSS.t31 VSS.t30 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X363 VOUT.t33 IBIAS.t104 a_n1962_4406.t2 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X364 a_3329_8823.t20 IBIAS.t105 a_3868_4185.t2 VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X365 VSS.t28 VSS.t26 a_3868_4185.t40 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X366 VDD.t45 VDD.t43 VDD.t45 VDD.t44 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X367 VDD.t42 VDD.t39 VDD.t41 VDD.t40 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X368 a_3868_4185.t1 IBIAS.t106 a_3329_8823.t31 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X369 a_3868_4185.t57 EN.t89 VSS.t222 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X370 a_3329_8823.t19 IBIAS.t107 a_3868_4185.t0 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X371 a_3868_4185.t56 EN.t90 VSS.t221 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X372 a_n1962_4406.t1 IBIAS.t108 VOUT.t27 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X373 VSS.t25 VSS.t24 a_n1962_4406.t60 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X374 VSS.t23 VSS.t21 VSS.t23 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X375 VSS.t220 EN.t91 a_8862_4192.t4 VSS.t216 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X376 a_n935_8875.t0 VN.t15 a_3329_8823.t44 VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X377 a_n1962_4406.t0 IBIAS.t109 VOUT.t59 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
R0 EN.n0 EN.t47 117.266
R1 EN.n3 EN.t69 117.266
R2 EN.n7 EN.t91 117.266
R3 EN.n11 EN.t85 117.266
R4 EN.n15 EN.t41 117.266
R5 EN.n38 EN.t38 117.266
R6 EN.n41 EN.t83 117.266
R7 EN.n44 EN.t25 117.266
R8 EN.n50 EN.t82 117.266
R9 EN.n56 EN.t24 117.266
R10 EN.n62 EN.t55 117.266
R11 EN.n68 EN.t1 117.266
R12 EN.n74 EN.t23 117.266
R13 EN.n80 EN.t73 117.266
R14 EN.n19 EN.t66 117.266
R15 EN.n22 EN.t72 117.266
R16 EN.n26 EN.t35 117.266
R17 EN.n30 EN.t39 117.266
R18 EN.n34 EN.t34 117.266
R19 EN.n87 EN.t58 117.266
R20 EN.n89 EN.t36 116.647
R21 EN.n88 EN.t31 116.647
R22 EN.n87 EN.t63 116.647
R23 EN.n2 EN.t19 116.647
R24 EN.n1 EN.t17 116.647
R25 EN.n0 EN.t50 116.647
R26 EN.n5 EN.t46 116.647
R27 EN.n4 EN.t44 116.647
R28 EN.n3 EN.t71 116.647
R29 EN.n9 EN.t65 116.647
R30 EN.n8 EN.t61 116.647
R31 EN.n7 EN.t0 116.647
R32 EN.n13 EN.t57 116.647
R33 EN.n12 EN.t56 116.647
R34 EN.n11 EN.t87 116.647
R35 EN.n17 EN.t10 116.647
R36 EN.n16 EN.t9 116.647
R37 EN.n15 EN.t45 116.647
R38 EN.n38 EN.t33 116.647
R39 EN.n39 EN.t84 116.647
R40 EN.n40 EN.t76 116.647
R41 EN.n41 EN.t60 116.647
R42 EN.n42 EN.t64 116.647
R43 EN.n43 EN.t51 116.647
R44 EN.n44 EN.t27 116.647
R45 EN.n45 EN.t30 116.647
R46 EN.n46 EN.t8 116.647
R47 EN.n47 EN.t68 116.647
R48 EN.n48 EN.t43 116.647
R49 EN.n50 EN.t59 116.647
R50 EN.n51 EN.t62 116.647
R51 EN.n52 EN.t49 116.647
R52 EN.n53 EN.t14 116.647
R53 EN.n54 EN.t12 116.647
R54 EN.n56 EN.t26 116.647
R55 EN.n57 EN.t29 116.647
R56 EN.n58 EN.t7 116.647
R57 EN.n59 EN.t67 116.647
R58 EN.n60 EN.t42 116.647
R59 EN.n62 EN.t28 116.647
R60 EN.n63 EN.t32 116.647
R61 EN.n64 EN.t18 116.647
R62 EN.n65 EN.t80 116.647
R63 EN.n66 EN.t75 116.647
R64 EN.n68 EN.t2 116.647
R65 EN.n69 EN.t3 116.647
R66 EN.n70 EN.t74 116.647
R67 EN.n71 EN.t40 116.647
R68 EN.n72 EN.t6 116.647
R69 EN.n74 EN.t4 116.647
R70 EN.n75 EN.t5 116.647
R71 EN.n76 EN.t88 116.647
R72 EN.n77 EN.t54 116.647
R73 EN.n78 EN.t52 116.647
R74 EN.n80 EN.t53 116.647
R75 EN.n81 EN.t11 116.647
R76 EN.n82 EN.t79 116.647
R77 EN.n19 EN.t21 116.647
R78 EN.n20 EN.t13 116.647
R79 EN.n21 EN.t48 116.647
R80 EN.n22 EN.t70 116.647
R81 EN.n23 EN.t22 116.647
R82 EN.n24 EN.t20 116.647
R83 EN.n26 EN.t90 116.647
R84 EN.n27 EN.t78 116.647
R85 EN.n28 EN.t16 116.647
R86 EN.n30 EN.t37 116.647
R87 EN.n31 EN.t86 116.647
R88 EN.n32 EN.t81 116.647
R89 EN.n34 EN.t89 116.647
R90 EN.n35 EN.t77 116.647
R91 EN.n36 EN.t15 116.647
R92 EN.n84 EN.n83 13.2346
R93 EN EN.n90 9.36508
R94 EN.n49 EN.n43 5.59733
R95 EN.n25 EN.n21 4.90021
R96 EN.n29 EN.n28 3.90565
R97 EN.n37 EN.n36 3.90565
R98 EN.n6 EN.n2 3.65983
R99 EN.n49 EN.n48 3.36238
R100 EN.n61 EN.n60 3.36238
R101 EN.n73 EN.n72 3.36238
R102 EN.n83 EN.n82 3.36238
R103 EN.n6 EN.n5 2.66526
R104 EN.n10 EN.n9 2.66526
R105 EN.n14 EN.n13 2.66526
R106 EN.n18 EN.n17 2.66526
R107 EN.n25 EN.n24 2.66526
R108 EN.n33 EN.n32 2.66526
R109 EN.n90 EN.n89 2.23017
R110 EN.n14 EN.n10 2.13093
R111 EN.n55 EN.n54 2.12199
R112 EN.n67 EN.n66 2.12199
R113 EN.n79 EN.n78 2.12199
R114 EN.n84 EN.n40 2.08834
R115 EN.n39 EN.n38 1.85887
R116 EN.n42 EN.n41 1.85887
R117 EN.n47 EN.n46 1.85887
R118 EN.n45 EN.n44 1.85887
R119 EN.n53 EN.n52 1.85887
R120 EN.n51 EN.n50 1.85887
R121 EN.n59 EN.n58 1.85887
R122 EN.n57 EN.n56 1.85887
R123 EN.n65 EN.n64 1.85887
R124 EN.n63 EN.n62 1.85887
R125 EN.n71 EN.n70 1.85887
R126 EN.n69 EN.n68 1.85887
R127 EN.n77 EN.n76 1.85887
R128 EN.n75 EN.n74 1.85887
R129 EN.n81 EN.n80 1.85887
R130 EN.n20 EN.n19 1.85887
R131 EN.n23 EN.n22 1.85887
R132 EN.n27 EN.n26 1.85887
R133 EN.n31 EN.n30 1.85887
R134 EN.n35 EN.n34 1.85887
R135 EN.n86 EN.n85 1.48383
R136 EN.n90 EN.n86 1.01147
R137 EN.n10 EN.n6 0.995065
R138 EN.n18 EN.n14 0.995065
R139 EN.n55 EN.n49 0.995065
R140 EN.n61 EN.n55 0.995065
R141 EN.n67 EN.n61 0.995065
R142 EN.n73 EN.n67 0.995065
R143 EN.n79 EN.n73 0.995065
R144 EN.n83 EN.n79 0.995065
R145 EN.n29 EN.n25 0.995065
R146 EN.n33 EN.n29 0.995065
R147 EN.n37 EN.n33 0.995065
R148 EN.n85 EN.n37 0.973326
R149 EN.n1 EN.n0 0.618487
R150 EN.n2 EN.n1 0.618487
R151 EN.n4 EN.n3 0.618487
R152 EN.n5 EN.n4 0.618487
R153 EN.n8 EN.n7 0.618487
R154 EN.n9 EN.n8 0.618487
R155 EN.n12 EN.n11 0.618487
R156 EN.n13 EN.n12 0.618487
R157 EN.n16 EN.n15 0.618487
R158 EN.n17 EN.n16 0.618487
R159 EN.n40 EN.n39 0.618487
R160 EN.n43 EN.n42 0.618487
R161 EN.n48 EN.n47 0.618487
R162 EN.n46 EN.n45 0.618487
R163 EN.n54 EN.n53 0.618487
R164 EN.n52 EN.n51 0.618487
R165 EN.n60 EN.n59 0.618487
R166 EN.n58 EN.n57 0.618487
R167 EN.n66 EN.n65 0.618487
R168 EN.n64 EN.n63 0.618487
R169 EN.n72 EN.n71 0.618487
R170 EN.n70 EN.n69 0.618487
R171 EN.n78 EN.n77 0.618487
R172 EN.n76 EN.n75 0.618487
R173 EN.n82 EN.n81 0.618487
R174 EN.n21 EN.n20 0.618487
R175 EN.n24 EN.n23 0.618487
R176 EN.n28 EN.n27 0.618487
R177 EN.n32 EN.n31 0.618487
R178 EN.n36 EN.n35 0.618487
R179 EN.n88 EN.n87 0.618487
R180 EN.n89 EN.n88 0.618487
R181 EN.n85 EN.n84 0.425821
R182 EN.n86 EN.n18 0.111913
R183 VSS.n1977 VSS.n1888 37142.3
R184 VSS.n2092 VSS.n1496 22163.5
R185 VSS.n2383 VSS.n123 1477.5
R186 VSS.n1376 VSS.n719 1419.56
R187 VSS.n1211 VSS.n825 1396.38
R188 VSS.n2192 VSS.n243 1384.79
R189 VSS.n2109 VSS.n668 1309.47
R190 VSS.n2129 VSS.n317 1303.68
R191 VSS.n661 VSS.n314 1303.68
R192 VSS.n2337 VSS.n165 1303.68
R193 VSS.n1494 VSS.n722 1303.68
R194 VSS.n1905 VSS.n1529 1263.12
R195 VSS.n187 VSS.n167 1245.74
R196 VSS.n2224 VSS.n213 1210.97
R197 VSS.n590 VSS.n211 1210.97
R198 VSS.n1207 VSS.n826 1210.97
R199 VSS.n2090 VSS.n1499 1187.79
R200 VSS.n1886 VSS.n1534 1158.82
R201 VSS.n1879 VSS.n1878 1158.82
R202 VSS.n1639 VSS.n127 1141.44
R203 VSS.n524 VSS.n523 788
R204 VSS.n568 VSS.n567 788
R205 VSS.n1663 VSS.n1662 788
R206 VSS.n1707 VSS.n1706 788
R207 VSS.n2335 VSS.n2226 712.073
R208 VSS.n165 VSS.n164 585
R209 VSS.n2333 VSS.n2332 585
R210 VSS.n2331 VSS.n2227 585
R211 VSS.n2335 VSS.n2227 585
R212 VSS.n2330 VSS.n2329 585
R213 VSS.n2328 VSS.n2327 585
R214 VSS.n2326 VSS.n2325 585
R215 VSS.n2324 VSS.n2323 585
R216 VSS.n2322 VSS.n2321 585
R217 VSS.n2320 VSS.n2319 585
R218 VSS.n2318 VSS.n2317 585
R219 VSS.n2316 VSS.n2315 585
R220 VSS.n2314 VSS.n2313 585
R221 VSS.n2312 VSS.n2311 585
R222 VSS.n2310 VSS.n2309 585
R223 VSS.n2308 VSS.n2307 585
R224 VSS.n2306 VSS.n2305 585
R225 VSS.n2304 VSS.n2303 585
R226 VSS.n2302 VSS.n2301 585
R227 VSS.n2300 VSS.n2299 585
R228 VSS.n2298 VSS.n2297 585
R229 VSS.n2296 VSS.n2295 585
R230 VSS.n2294 VSS.n2293 585
R231 VSS.n2292 VSS.n2291 585
R232 VSS.n2290 VSS.n2289 585
R233 VSS.n2288 VSS.n2287 585
R234 VSS.n2286 VSS.n2285 585
R235 VSS.n2284 VSS.n2283 585
R236 VSS.n2282 VSS.n2281 585
R237 VSS.n2280 VSS.n2279 585
R238 VSS.n2278 VSS.n2277 585
R239 VSS.n2276 VSS.n2275 585
R240 VSS.n2274 VSS.n2273 585
R241 VSS.n2272 VSS.n2271 585
R242 VSS.n2270 VSS.n2269 585
R243 VSS.n2268 VSS.n2267 585
R244 VSS.n2266 VSS.n2265 585
R245 VSS.n2264 VSS.n2263 585
R246 VSS.n2262 VSS.n2261 585
R247 VSS.n2260 VSS.n2259 585
R248 VSS.n2258 VSS.n2257 585
R249 VSS.n2256 VSS.n2255 585
R250 VSS.n2254 VSS.n187 585
R251 VSS.n2335 VSS.n187 585
R252 VSS.n2253 VSS.n167 585
R253 VSS.n2336 VSS.n167 585
R254 VSS.n2252 VSS.n2251 585
R255 VSS.n2251 VSS.n166 585
R256 VSS.n2250 VSS.n162 585
R257 VSS.n2342 VSS.n162 585
R258 VSS.n2249 VSS.n161 585
R259 VSS.n2343 VSS.n161 585
R260 VSS.n2248 VSS.n160 585
R261 VSS.n2344 VSS.n160 585
R262 VSS.n2247 VSS.n2246 585
R263 VSS.n2246 VSS.n159 585
R264 VSS.n2245 VSS.n155 585
R265 VSS.n2350 VSS.n155 585
R266 VSS.n2244 VSS.n154 585
R267 VSS.n2351 VSS.n154 585
R268 VSS.n2243 VSS.n153 585
R269 VSS.n2352 VSS.n153 585
R270 VSS.n2242 VSS.n2241 585
R271 VSS.n2241 VSS.n152 585
R272 VSS.n2240 VSS.n148 585
R273 VSS.n2358 VSS.n148 585
R274 VSS.n2239 VSS.n147 585
R275 VSS.n2359 VSS.n147 585
R276 VSS.n2238 VSS.n146 585
R277 VSS.n2360 VSS.n146 585
R278 VSS.n2237 VSS.n2236 585
R279 VSS.n2236 VSS.n145 585
R280 VSS.n2235 VSS.n141 585
R281 VSS.n2366 VSS.n141 585
R282 VSS.n2234 VSS.n140 585
R283 VSS.n2367 VSS.n140 585
R284 VSS.n2233 VSS.n139 585
R285 VSS.n2368 VSS.n139 585
R286 VSS.n2232 VSS.n2231 585
R287 VSS.n2231 VSS.n135 585
R288 VSS.n2230 VSS.n134 585
R289 VSS.n2374 VSS.n134 585
R290 VSS.n2229 VSS.n133 585
R291 VSS.n2375 VSS.n133 585
R292 VSS.n2228 VSS.n132 585
R293 VSS.n2376 VSS.n132 585
R294 VSS.n124 VSS.n122 585
R295 VSS.n126 VSS.n124 585
R296 VSS.n2384 VSS.n2383 585
R297 VSS.n2383 VSS.n2382 585
R298 VSS.n123 VSS.n121 585
R299 VSS.n1715 VSS.n1714 585
R300 VSS.n1713 VSS.n1638 585
R301 VSS.n1712 VSS.n1711 585
R302 VSS.n1710 VSS.n1709 585
R303 VSS.n1708 VSS.n1707 585
R304 VSS.n1706 VSS.n1705 585
R305 VSS.n1704 VSS.n1703 585
R306 VSS.n1702 VSS.n1701 585
R307 VSS.n1700 VSS.n1699 585
R308 VSS.n1698 VSS.n1697 585
R309 VSS.n1696 VSS.n1695 585
R310 VSS.n1694 VSS.n1693 585
R311 VSS.n1692 VSS.n1691 585
R312 VSS.n1690 VSS.n1689 585
R313 VSS.n1688 VSS.n1687 585
R314 VSS.n1686 VSS.n1685 585
R315 VSS.n1684 VSS.n1683 585
R316 VSS.n1682 VSS.n1681 585
R317 VSS.n1680 VSS.n1679 585
R318 VSS.n1678 VSS.n1677 585
R319 VSS.n1676 VSS.n1675 585
R320 VSS.n1674 VSS.n1673 585
R321 VSS.n1672 VSS.n1671 585
R322 VSS.n1670 VSS.n1669 585
R323 VSS.n1668 VSS.n1667 585
R324 VSS.n1666 VSS.n1665 585
R325 VSS.n1664 VSS.n1663 585
R326 VSS.n1662 VSS.n1661 585
R327 VSS.n1660 VSS.n1659 585
R328 VSS.n1658 VSS.n1657 585
R329 VSS.n1656 VSS.n1655 585
R330 VSS.n1654 VSS.n1653 585
R331 VSS.n1652 VSS.n1651 585
R332 VSS.n1650 VSS.n1649 585
R333 VSS.n1648 VSS.n1647 585
R334 VSS.n1646 VSS.n1645 585
R335 VSS.n1644 VSS.n1643 585
R336 VSS.n1642 VSS.n1641 585
R337 VSS.n1640 VSS.n1639 585
R338 VSS.n129 VSS.n127 585
R339 VSS.n1718 VSS.n127 585
R340 VSS.n2381 VSS.n2380 585
R341 VSS.n2382 VSS.n2381 585
R342 VSS.n2379 VSS.n128 585
R343 VSS.n128 VSS.n126 585
R344 VSS.n2378 VSS.n2377 585
R345 VSS.n2377 VSS.n2376 585
R346 VSS.n131 VSS.n130 585
R347 VSS.n2375 VSS.n131 585
R348 VSS.n2373 VSS.n2372 585
R349 VSS.n2374 VSS.n2373 585
R350 VSS.n2371 VSS.n136 585
R351 VSS.n136 VSS.n135 585
R352 VSS.n2370 VSS.n2369 585
R353 VSS.n2369 VSS.n2368 585
R354 VSS.n138 VSS.n137 585
R355 VSS.n2367 VSS.n138 585
R356 VSS.n2365 VSS.n2364 585
R357 VSS.n2366 VSS.n2365 585
R358 VSS.n2363 VSS.n142 585
R359 VSS.n145 VSS.n142 585
R360 VSS.n2362 VSS.n2361 585
R361 VSS.n2361 VSS.n2360 585
R362 VSS.n144 VSS.n143 585
R363 VSS.n2359 VSS.n144 585
R364 VSS.n2357 VSS.n2356 585
R365 VSS.n2358 VSS.n2357 585
R366 VSS.n2355 VSS.n149 585
R367 VSS.n152 VSS.n149 585
R368 VSS.n2354 VSS.n2353 585
R369 VSS.n2353 VSS.n2352 585
R370 VSS.n151 VSS.n150 585
R371 VSS.n2351 VSS.n151 585
R372 VSS.n2349 VSS.n2348 585
R373 VSS.n2350 VSS.n2349 585
R374 VSS.n2347 VSS.n156 585
R375 VSS.n159 VSS.n156 585
R376 VSS.n2346 VSS.n2345 585
R377 VSS.n2345 VSS.n2344 585
R378 VSS.n158 VSS.n157 585
R379 VSS.n2343 VSS.n158 585
R380 VSS.n2341 VSS.n2340 585
R381 VSS.n2342 VSS.n2341 585
R382 VSS.n2339 VSS.n163 585
R383 VSS.n166 VSS.n163 585
R384 VSS.n2338 VSS.n2337 585
R385 VSS.n2337 VSS.n2336 585
R386 VSS.n1785 VSS.n1617 585
R387 VSS.n1617 VSS.n1616 585
R388 VSS.n1784 VSS.n1783 585
R389 VSS.n1783 VSS.n1782 585
R390 VSS.n1779 VSS.n1778 585
R391 VSS.n1780 VSS.n1779 585
R392 VSS.n1777 VSS.n1720 585
R393 VSS.n1720 VSS.n1719 585
R394 VSS.n1776 VSS.n1775 585
R395 VSS.n1775 VSS.n125 585
R396 VSS.n1878 VSS.n1536 585
R397 VSS.n1878 VSS.n1531 585
R398 VSS.n1877 VSS.n1538 585
R399 VSS.n1877 VSS.n1876 585
R400 VSS.n1721 VSS.n1537 585
R401 VSS.n1539 VSS.n1537 585
R402 VSS.n1722 VSS.n1543 585
R403 VSS.n1870 VSS.n1543 585
R404 VSS.n1723 VSS.n1544 585
R405 VSS.n1869 VSS.n1544 585
R406 VSS.n1724 VSS.n1545 585
R407 VSS.n1868 VSS.n1545 585
R408 VSS.n1726 VSS.n1725 585
R409 VSS.n1725 VSS.n1546 585
R410 VSS.n1727 VSS.n1550 585
R411 VSS.n1862 VSS.n1550 585
R412 VSS.n1728 VSS.n1551 585
R413 VSS.n1861 VSS.n1551 585
R414 VSS.n1729 VSS.n1552 585
R415 VSS.n1860 VSS.n1552 585
R416 VSS.n1731 VSS.n1730 585
R417 VSS.n1730 VSS.n1553 585
R418 VSS.n1732 VSS.n1557 585
R419 VSS.n1854 VSS.n1557 585
R420 VSS.n1733 VSS.n1558 585
R421 VSS.n1853 VSS.n1558 585
R422 VSS.n1734 VSS.n1559 585
R423 VSS.n1852 VSS.n1559 585
R424 VSS.n1736 VSS.n1735 585
R425 VSS.n1735 VSS.n1560 585
R426 VSS.n1737 VSS.n1564 585
R427 VSS.n1846 VSS.n1564 585
R428 VSS.n1738 VSS.n1565 585
R429 VSS.n1845 VSS.n1565 585
R430 VSS.n1739 VSS.n1566 585
R431 VSS.n1844 VSS.n1566 585
R432 VSS.n1741 VSS.n1740 585
R433 VSS.n1740 VSS.n1567 585
R434 VSS.n1742 VSS.n1571 585
R435 VSS.n1838 VSS.n1571 585
R436 VSS.n1743 VSS.n1572 585
R437 VSS.n1837 VSS.n1572 585
R438 VSS.n1744 VSS.n1573 585
R439 VSS.n1836 VSS.n1573 585
R440 VSS.n1746 VSS.n1745 585
R441 VSS.n1745 VSS.n1574 585
R442 VSS.n1747 VSS.n1578 585
R443 VSS.n1830 VSS.n1578 585
R444 VSS.n1748 VSS.n1579 585
R445 VSS.n1829 VSS.n1579 585
R446 VSS.n1749 VSS.n1580 585
R447 VSS.n1828 VSS.n1580 585
R448 VSS.n1751 VSS.n1750 585
R449 VSS.n1750 VSS.n1581 585
R450 VSS.n1752 VSS.n1585 585
R451 VSS.n1822 VSS.n1585 585
R452 VSS.n1753 VSS.n1586 585
R453 VSS.n1821 VSS.n1586 585
R454 VSS.n1754 VSS.n1587 585
R455 VSS.n1820 VSS.n1587 585
R456 VSS.n1756 VSS.n1755 585
R457 VSS.n1755 VSS.n1588 585
R458 VSS.n1757 VSS.n1592 585
R459 VSS.n1814 VSS.n1592 585
R460 VSS.n1758 VSS.n1593 585
R461 VSS.n1813 VSS.n1593 585
R462 VSS.n1759 VSS.n1594 585
R463 VSS.n1812 VSS.n1594 585
R464 VSS.n1761 VSS.n1760 585
R465 VSS.n1760 VSS.n1595 585
R466 VSS.n1762 VSS.n1599 585
R467 VSS.n1806 VSS.n1599 585
R468 VSS.n1763 VSS.n1600 585
R469 VSS.n1805 VSS.n1600 585
R470 VSS.n1764 VSS.n1601 585
R471 VSS.n1804 VSS.n1601 585
R472 VSS.n1766 VSS.n1765 585
R473 VSS.n1765 VSS.n1602 585
R474 VSS.n1767 VSS.n1606 585
R475 VSS.n1798 VSS.n1606 585
R476 VSS.n1768 VSS.n1607 585
R477 VSS.n1797 VSS.n1607 585
R478 VSS.n1769 VSS.n1608 585
R479 VSS.n1796 VSS.n1608 585
R480 VSS.n1771 VSS.n1770 585
R481 VSS.n1770 VSS.n1609 585
R482 VSS.n1772 VSS.n1613 585
R483 VSS.n1790 VSS.n1613 585
R484 VSS.n1773 VSS.n1614 585
R485 VSS.n1789 VSS.n1614 585
R486 VSS.n1774 VSS.n1615 585
R487 VSS.n1788 VSS.n1615 585
R488 VSS.n1787 VSS.n1786 585
R489 VSS.n1788 VSS.n1787 585
R490 VSS.n1612 VSS.n1611 585
R491 VSS.n1789 VSS.n1612 585
R492 VSS.n1792 VSS.n1791 585
R493 VSS.n1791 VSS.n1790 585
R494 VSS.n1793 VSS.n1610 585
R495 VSS.n1610 VSS.n1609 585
R496 VSS.n1795 VSS.n1794 585
R497 VSS.n1796 VSS.n1795 585
R498 VSS.n1605 VSS.n1604 585
R499 VSS.n1797 VSS.n1605 585
R500 VSS.n1800 VSS.n1799 585
R501 VSS.n1799 VSS.n1798 585
R502 VSS.n1801 VSS.n1603 585
R503 VSS.n1603 VSS.n1602 585
R504 VSS.n1803 VSS.n1802 585
R505 VSS.n1804 VSS.n1803 585
R506 VSS.n1598 VSS.n1597 585
R507 VSS.n1805 VSS.n1598 585
R508 VSS.n1808 VSS.n1807 585
R509 VSS.n1807 VSS.n1806 585
R510 VSS.n1809 VSS.n1596 585
R511 VSS.n1596 VSS.n1595 585
R512 VSS.n1811 VSS.n1810 585
R513 VSS.n1812 VSS.n1811 585
R514 VSS.n1591 VSS.n1590 585
R515 VSS.n1813 VSS.n1591 585
R516 VSS.n1816 VSS.n1815 585
R517 VSS.n1815 VSS.n1814 585
R518 VSS.n1817 VSS.n1589 585
R519 VSS.n1589 VSS.n1588 585
R520 VSS.n1819 VSS.n1818 585
R521 VSS.n1820 VSS.n1819 585
R522 VSS.n1584 VSS.n1583 585
R523 VSS.n1821 VSS.n1584 585
R524 VSS.n1824 VSS.n1823 585
R525 VSS.n1823 VSS.n1822 585
R526 VSS.n1825 VSS.n1582 585
R527 VSS.n1582 VSS.n1581 585
R528 VSS.n1827 VSS.n1826 585
R529 VSS.n1828 VSS.n1827 585
R530 VSS.n1577 VSS.n1576 585
R531 VSS.n1829 VSS.n1577 585
R532 VSS.n1832 VSS.n1831 585
R533 VSS.n1831 VSS.n1830 585
R534 VSS.n1833 VSS.n1575 585
R535 VSS.n1575 VSS.n1574 585
R536 VSS.n1835 VSS.n1834 585
R537 VSS.n1836 VSS.n1835 585
R538 VSS.n1570 VSS.n1569 585
R539 VSS.n1837 VSS.n1570 585
R540 VSS.n1840 VSS.n1839 585
R541 VSS.n1839 VSS.n1838 585
R542 VSS.n1841 VSS.n1568 585
R543 VSS.n1568 VSS.n1567 585
R544 VSS.n1843 VSS.n1842 585
R545 VSS.n1844 VSS.n1843 585
R546 VSS.n1563 VSS.n1562 585
R547 VSS.n1845 VSS.n1563 585
R548 VSS.n1848 VSS.n1847 585
R549 VSS.n1847 VSS.n1846 585
R550 VSS.n1849 VSS.n1561 585
R551 VSS.n1561 VSS.n1560 585
R552 VSS.n1851 VSS.n1850 585
R553 VSS.n1852 VSS.n1851 585
R554 VSS.n1556 VSS.n1555 585
R555 VSS.n1853 VSS.n1556 585
R556 VSS.n1856 VSS.n1855 585
R557 VSS.n1855 VSS.n1854 585
R558 VSS.n1857 VSS.n1554 585
R559 VSS.n1554 VSS.n1553 585
R560 VSS.n1859 VSS.n1858 585
R561 VSS.n1860 VSS.n1859 585
R562 VSS.n1549 VSS.n1548 585
R563 VSS.n1861 VSS.n1549 585
R564 VSS.n1864 VSS.n1863 585
R565 VSS.n1863 VSS.n1862 585
R566 VSS.n1865 VSS.n1547 585
R567 VSS.n1547 VSS.n1546 585
R568 VSS.n1867 VSS.n1866 585
R569 VSS.n1868 VSS.n1867 585
R570 VSS.n1542 VSS.n1541 585
R571 VSS.n1869 VSS.n1542 585
R572 VSS.n1872 VSS.n1871 585
R573 VSS.n1871 VSS.n1870 585
R574 VSS.n1873 VSS.n1540 585
R575 VSS.n1540 VSS.n1539 585
R576 VSS.n1875 VSS.n1874 585
R577 VSS.n1876 VSS.n1875 585
R578 VSS.n1535 VSS.n1534 585
R579 VSS.n1534 VSS.n1531 585
R580 VSS.n1886 VSS.n1885 585
R581 VSS.n1884 VSS.n1533 585
R582 VSS.n1883 VSS.n1532 585
R583 VSS.n1888 VSS.n1532 585
R584 VSS.n1882 VSS.n1881 585
R585 VSS.n1880 VSS.n1879 585
R586 VSS.n2090 VSS.n2089 585
R587 VSS.n2088 VSS.n1498 585
R588 VSS.n2087 VSS.n1497 585
R589 VSS.n2092 VSS.n1497 585
R590 VSS.n2086 VSS.n2085 585
R591 VSS.n2084 VSS.n2083 585
R592 VSS.n2082 VSS.n2081 585
R593 VSS.n2080 VSS.n2079 585
R594 VSS.n2078 VSS.n2077 585
R595 VSS.n2076 VSS.n2075 585
R596 VSS.n2074 VSS.n2073 585
R597 VSS.n2072 VSS.n2071 585
R598 VSS.n2070 VSS.n2069 585
R599 VSS.n2068 VSS.n2067 585
R600 VSS.n2066 VSS.n2065 585
R601 VSS.n2064 VSS.n2063 585
R602 VSS.n2062 VSS.n2061 585
R603 VSS.n2060 VSS.n2059 585
R604 VSS.n2058 VSS.n2057 585
R605 VSS.n2056 VSS.n2055 585
R606 VSS.n2054 VSS.n2053 585
R607 VSS.n2052 VSS.n2051 585
R608 VSS.n2050 VSS.n2049 585
R609 VSS.n2048 VSS.n2047 585
R610 VSS.n2046 VSS.n2045 585
R611 VSS.n2044 VSS.n2043 585
R612 VSS.n2042 VSS.n2041 585
R613 VSS.n2040 VSS.n2039 585
R614 VSS.n676 VSS.n675 585
R615 VSS.n2095 VSS.n2094 585
R616 VSS.n2096 VSS.n674 585
R617 VSS.n2092 VSS.n674 585
R618 VSS.n1975 VSS.n1974 585
R619 VSS.n1961 VSS.n1903 585
R620 VSS.n1960 VSS.n1959 585
R621 VSS.n1958 VSS.n1957 585
R622 VSS.n1956 VSS.n1955 585
R623 VSS.n1954 VSS.n1953 585
R624 VSS.n1952 VSS.n1951 585
R625 VSS.n1950 VSS.n1949 585
R626 VSS.n1948 VSS.n1947 585
R627 VSS.n1946 VSS.n1945 585
R628 VSS.n1944 VSS.n1943 585
R629 VSS.n1942 VSS.n1941 585
R630 VSS.n1940 VSS.n1939 585
R631 VSS.n1938 VSS.n1937 585
R632 VSS.n1936 VSS.n1935 585
R633 VSS.n1934 VSS.n1933 585
R634 VSS.n1932 VSS.n1931 585
R635 VSS.n1930 VSS.n1929 585
R636 VSS.n1928 VSS.n1927 585
R637 VSS.n1926 VSS.n1925 585
R638 VSS.n1924 VSS.n1923 585
R639 VSS.n1922 VSS.n1921 585
R640 VSS.n1920 VSS.n1919 585
R641 VSS.n1918 VSS.n1917 585
R642 VSS.n1916 VSS.n1915 585
R643 VSS.n1914 VSS.n1913 585
R644 VSS.n1912 VSS.n1911 585
R645 VSS.n1910 VSS.n1909 585
R646 VSS.n1908 VSS.n1907 585
R647 VSS.n1906 VSS.n1905 585
R648 VSS.n1529 VSS.n1528 585
R649 VSS.n1978 VSS.n1529 585
R650 VSS.n1981 VSS.n1980 585
R651 VSS.n1980 VSS.n1979 585
R652 VSS.n1982 VSS.n1527 585
R653 VSS.n1527 VSS.n1526 585
R654 VSS.n1984 VSS.n1983 585
R655 VSS.n1985 VSS.n1984 585
R656 VSS.n1525 VSS.n1524 585
R657 VSS.n1986 VSS.n1525 585
R658 VSS.n1989 VSS.n1988 585
R659 VSS.n1988 VSS.n1987 585
R660 VSS.n1990 VSS.n1523 585
R661 VSS.n1523 VSS.n1522 585
R662 VSS.n1992 VSS.n1991 585
R663 VSS.n1993 VSS.n1992 585
R664 VSS.n1521 VSS.n1520 585
R665 VSS.n1994 VSS.n1521 585
R666 VSS.n1997 VSS.n1996 585
R667 VSS.n1996 VSS.n1995 585
R668 VSS.n1998 VSS.n1519 585
R669 VSS.n1519 VSS.n1518 585
R670 VSS.n2000 VSS.n1999 585
R671 VSS.n2001 VSS.n2000 585
R672 VSS.n1517 VSS.n1516 585
R673 VSS.n2002 VSS.n1517 585
R674 VSS.n2005 VSS.n2004 585
R675 VSS.n2004 VSS.n2003 585
R676 VSS.n2006 VSS.n1515 585
R677 VSS.n1515 VSS.n1514 585
R678 VSS.n2008 VSS.n2007 585
R679 VSS.n2009 VSS.n2008 585
R680 VSS.n1513 VSS.n1512 585
R681 VSS.n2010 VSS.n1513 585
R682 VSS.n2013 VSS.n2012 585
R683 VSS.n2012 VSS.n2011 585
R684 VSS.n2014 VSS.n1511 585
R685 VSS.n1511 VSS.n1510 585
R686 VSS.n2016 VSS.n2015 585
R687 VSS.n2017 VSS.n2016 585
R688 VSS.n1509 VSS.n1508 585
R689 VSS.n2018 VSS.n1509 585
R690 VSS.n2021 VSS.n2020 585
R691 VSS.n2020 VSS.n2019 585
R692 VSS.n2022 VSS.n1507 585
R693 VSS.n1507 VSS.n1506 585
R694 VSS.n2024 VSS.n2023 585
R695 VSS.n2025 VSS.n2024 585
R696 VSS.n1505 VSS.n1504 585
R697 VSS.n2026 VSS.n1505 585
R698 VSS.n2029 VSS.n2028 585
R699 VSS.n2028 VSS.n2027 585
R700 VSS.n2030 VSS.n1503 585
R701 VSS.n1503 VSS.n1502 585
R702 VSS.n2032 VSS.n2031 585
R703 VSS.n2033 VSS.n2032 585
R704 VSS.n1501 VSS.n1500 585
R705 VSS.n2034 VSS.n1501 585
R706 VSS.n2037 VSS.n2036 585
R707 VSS.n2036 VSS.n2035 585
R708 VSS.n2038 VSS.n1499 585
R709 VSS.n1499 VSS.n677 585
R710 VSS.n2127 VSS.n317 585
R711 VSS.n2126 VSS.n2125 585
R712 VSS.n320 VSS.n319 585
R713 VSS.n2123 VSS.n320 585
R714 VSS.n345 VSS.n344 585
R715 VSS.n347 VSS.n346 585
R716 VSS.n349 VSS.n348 585
R717 VSS.n351 VSS.n350 585
R718 VSS.n353 VSS.n352 585
R719 VSS.n355 VSS.n354 585
R720 VSS.n357 VSS.n356 585
R721 VSS.n359 VSS.n358 585
R722 VSS.n361 VSS.n360 585
R723 VSS.n363 VSS.n362 585
R724 VSS.n365 VSS.n364 585
R725 VSS.n367 VSS.n366 585
R726 VSS.n369 VSS.n368 585
R727 VSS.n371 VSS.n370 585
R728 VSS.n373 VSS.n372 585
R729 VSS.n375 VSS.n374 585
R730 VSS.n377 VSS.n376 585
R731 VSS.n379 VSS.n378 585
R732 VSS.n381 VSS.n380 585
R733 VSS.n383 VSS.n382 585
R734 VSS.n385 VSS.n384 585
R735 VSS.n387 VSS.n386 585
R736 VSS.n389 VSS.n388 585
R737 VSS.n391 VSS.n390 585
R738 VSS.n393 VSS.n392 585
R739 VSS.n395 VSS.n394 585
R740 VSS.n397 VSS.n396 585
R741 VSS.n399 VSS.n398 585
R742 VSS.n401 VSS.n400 585
R743 VSS.n403 VSS.n402 585
R744 VSS.n405 VSS.n404 585
R745 VSS.n407 VSS.n406 585
R746 VSS.n409 VSS.n408 585
R747 VSS.n411 VSS.n410 585
R748 VSS.n413 VSS.n412 585
R749 VSS.n415 VSS.n414 585
R750 VSS.n417 VSS.n416 585
R751 VSS.n419 VSS.n418 585
R752 VSS.n421 VSS.n420 585
R753 VSS.n423 VSS.n422 585
R754 VSS.n425 VSS.n424 585
R755 VSS.n427 VSS.n426 585
R756 VSS.n429 VSS.n428 585
R757 VSS.n430 VSS.n343 585
R758 VSS.n661 VSS.n660 585
R759 VSS.n2123 VSS.n661 585
R760 VSS.n659 VSS.n314 585
R761 VSS.n2130 VSS.n314 585
R762 VSS.n658 VSS.n657 585
R763 VSS.n657 VSS.n656 585
R764 VSS.n654 VSS.n653 585
R765 VSS.n654 VSS.n307 585
R766 VSS.n652 VSS.n306 585
R767 VSS.n2138 VSS.n306 585
R768 VSS.n651 VSS.n650 585
R769 VSS.n650 VSS.n649 585
R770 VSS.n648 VSS.n298 585
R771 VSS.n2144 VSS.n298 585
R772 VSS.n647 VSS.n646 585
R773 VSS.n646 VSS.n645 585
R774 VSS.n643 VSS.n642 585
R775 VSS.n643 VSS.n292 585
R776 VSS.n641 VSS.n291 585
R777 VSS.n2152 VSS.n291 585
R778 VSS.n640 VSS.n639 585
R779 VSS.n639 VSS.n638 585
R780 VSS.n636 VSS.n284 585
R781 VSS.n2158 VSS.n284 585
R782 VSS.n635 VSS.n634 585
R783 VSS.n634 VSS.n283 585
R784 VSS.n633 VSS.n632 585
R785 VSS.n633 VSS.n276 585
R786 VSS.n631 VSS.n275 585
R787 VSS.n2166 VSS.n275 585
R788 VSS.n630 VSS.n629 585
R789 VSS.n629 VSS.n628 585
R790 VSS.n627 VSS.n267 585
R791 VSS.n2172 VSS.n267 585
R792 VSS.n626 VSS.n625 585
R793 VSS.n625 VSS.n266 585
R794 VSS.n624 VSS.n623 585
R795 VSS.n624 VSS.n259 585
R796 VSS.n622 VSS.n258 585
R797 VSS.n2180 VSS.n258 585
R798 VSS.n621 VSS.n620 585
R799 VSS.n620 VSS.n619 585
R800 VSS.n618 VSS.n248 585
R801 VSS.n2186 VSS.n248 585
R802 VSS.n617 VSS.n616 585
R803 VSS.n616 VSS.n615 585
R804 VSS.n613 VSS.n612 585
R805 VSS.n613 VSS.n242 585
R806 VSS.n611 VSS.n241 585
R807 VSS.n2194 VSS.n241 585
R808 VSS.n610 VSS.n240 585
R809 VSS.n2195 VSS.n240 585
R810 VSS.n609 VSS.n608 585
R811 VSS.n608 VSS.n235 585
R812 VSS.n607 VSS.n234 585
R813 VSS.n2201 VSS.n234 585
R814 VSS.n606 VSS.n233 585
R815 VSS.n2202 VSS.n233 585
R816 VSS.n605 VSS.n232 585
R817 VSS.n2203 VSS.n232 585
R818 VSS.n604 VSS.n603 585
R819 VSS.n603 VSS.n228 585
R820 VSS.n602 VSS.n227 585
R821 VSS.n2209 VSS.n227 585
R822 VSS.n601 VSS.n226 585
R823 VSS.n2210 VSS.n226 585
R824 VSS.n600 VSS.n225 585
R825 VSS.n2211 VSS.n225 585
R826 VSS.n599 VSS.n598 585
R827 VSS.n598 VSS.n221 585
R828 VSS.n597 VSS.n220 585
R829 VSS.n2217 VSS.n220 585
R830 VSS.n596 VSS.n219 585
R831 VSS.n2218 VSS.n219 585
R832 VSS.n595 VSS.n218 585
R833 VSS.n2219 VSS.n218 585
R834 VSS.n594 VSS.n593 585
R835 VSS.n593 VSS.n212 585
R836 VSS.n592 VSS.n211 585
R837 VSS.n2225 VSS.n211 585
R838 VSS.n591 VSS.n590 585
R839 VSS.n589 VSS.n588 585
R840 VSS.n587 VSS.n586 585
R841 VSS.n585 VSS.n584 585
R842 VSS.n583 VSS.n582 585
R843 VSS.n581 VSS.n580 585
R844 VSS.n579 VSS.n578 585
R845 VSS.n577 VSS.n576 585
R846 VSS.n575 VSS.n574 585
R847 VSS.n573 VSS.n572 585
R848 VSS.n571 VSS.n570 585
R849 VSS.n569 VSS.n568 585
R850 VSS.n567 VSS.n566 585
R851 VSS.n565 VSS.n564 585
R852 VSS.n563 VSS.n562 585
R853 VSS.n561 VSS.n560 585
R854 VSS.n559 VSS.n558 585
R855 VSS.n557 VSS.n556 585
R856 VSS.n555 VSS.n554 585
R857 VSS.n553 VSS.n552 585
R858 VSS.n551 VSS.n550 585
R859 VSS.n549 VSS.n548 585
R860 VSS.n547 VSS.n546 585
R861 VSS.n545 VSS.n544 585
R862 VSS.n543 VSS.n542 585
R863 VSS.n541 VSS.n540 585
R864 VSS.n539 VSS.n538 585
R865 VSS.n537 VSS.n536 585
R866 VSS.n535 VSS.n534 585
R867 VSS.n533 VSS.n532 585
R868 VSS.n531 VSS.n530 585
R869 VSS.n529 VSS.n528 585
R870 VSS.n527 VSS.n526 585
R871 VSS.n525 VSS.n524 585
R872 VSS.n523 VSS.n522 585
R873 VSS.n521 VSS.n520 585
R874 VSS.n519 VSS.n518 585
R875 VSS.n517 VSS.n516 585
R876 VSS.n515 VSS.n514 585
R877 VSS.n513 VSS.n512 585
R878 VSS.n511 VSS.n510 585
R879 VSS.n509 VSS.n508 585
R880 VSS.n507 VSS.n506 585
R881 VSS.n505 VSS.n504 585
R882 VSS.n503 VSS.n502 585
R883 VSS.n215 VSS.n213 585
R884 VSS.n2224 VSS.n2223 585
R885 VSS.n2225 VSS.n2224 585
R886 VSS.n2222 VSS.n214 585
R887 VSS.n214 VSS.n212 585
R888 VSS.n2221 VSS.n2220 585
R889 VSS.n2220 VSS.n2219 585
R890 VSS.n217 VSS.n216 585
R891 VSS.n2218 VSS.n217 585
R892 VSS.n2216 VSS.n2215 585
R893 VSS.n2217 VSS.n2216 585
R894 VSS.n2214 VSS.n222 585
R895 VSS.n222 VSS.n221 585
R896 VSS.n2213 VSS.n2212 585
R897 VSS.n2212 VSS.n2211 585
R898 VSS.n224 VSS.n223 585
R899 VSS.n2210 VSS.n224 585
R900 VSS.n2208 VSS.n2207 585
R901 VSS.n2209 VSS.n2208 585
R902 VSS.n2206 VSS.n229 585
R903 VSS.n229 VSS.n228 585
R904 VSS.n2205 VSS.n2204 585
R905 VSS.n2204 VSS.n2203 585
R906 VSS.n231 VSS.n230 585
R907 VSS.n2202 VSS.n231 585
R908 VSS.n2200 VSS.n2199 585
R909 VSS.n2201 VSS.n2200 585
R910 VSS.n2198 VSS.n236 585
R911 VSS.n236 VSS.n235 585
R912 VSS.n2197 VSS.n2196 585
R913 VSS.n2196 VSS.n2195 585
R914 VSS.n238 VSS.n237 585
R915 VSS.n2194 VSS.n238 585
R916 VSS.n253 VSS.n252 585
R917 VSS.n252 VSS.n242 585
R918 VSS.n254 VSS.n250 585
R919 VSS.n615 VSS.n250 585
R920 VSS.n2185 VSS.n2184 585
R921 VSS.n2186 VSS.n2185 585
R922 VSS.n2183 VSS.n251 585
R923 VSS.n619 VSS.n251 585
R924 VSS.n2182 VSS.n2181 585
R925 VSS.n2181 VSS.n2180 585
R926 VSS.n256 VSS.n255 585
R927 VSS.n259 VSS.n256 585
R928 VSS.n271 VSS.n269 585
R929 VSS.n269 VSS.n266 585
R930 VSS.n2171 VSS.n2170 585
R931 VSS.n2172 VSS.n2171 585
R932 VSS.n2169 VSS.n270 585
R933 VSS.n628 VSS.n270 585
R934 VSS.n2168 VSS.n2167 585
R935 VSS.n2167 VSS.n2166 585
R936 VSS.n273 VSS.n272 585
R937 VSS.n276 VSS.n273 585
R938 VSS.n287 VSS.n285 585
R939 VSS.n285 VSS.n283 585
R940 VSS.n2157 VSS.n2156 585
R941 VSS.n2158 VSS.n2157 585
R942 VSS.n2155 VSS.n286 585
R943 VSS.n638 VSS.n286 585
R944 VSS.n2154 VSS.n2153 585
R945 VSS.n2153 VSS.n2152 585
R946 VSS.n289 VSS.n288 585
R947 VSS.n292 VSS.n289 585
R948 VSS.n302 VSS.n300 585
R949 VSS.n645 VSS.n300 585
R950 VSS.n2143 VSS.n2142 585
R951 VSS.n2144 VSS.n2143 585
R952 VSS.n2141 VSS.n301 585
R953 VSS.n649 VSS.n301 585
R954 VSS.n2140 VSS.n2139 585
R955 VSS.n2139 VSS.n2138 585
R956 VSS.n304 VSS.n303 585
R957 VSS.n307 VSS.n304 585
R958 VSS.n318 VSS.n316 585
R959 VSS.n656 VSS.n316 585
R960 VSS.n2129 VSS.n2128 585
R961 VSS.n2130 VSS.n2129 585
R962 VSS.n2105 VSS.n2104 585
R963 VSS.n2103 VSS.n673 585
R964 VSS.n2102 VSS.n672 585
R965 VSS.n2107 VSS.n672 585
R966 VSS.n2101 VSS.n2100 585
R967 VSS.n2099 VSS.n2098 585
R968 VSS.n2097 VSS.n668 585
R969 VSS.n2107 VSS.n668 585
R970 VSS.n2110 VSS.n2109 585
R971 VSS.n2109 VSS.n2108 585
R972 VSS.n2111 VSS.n666 585
R973 VSS.n669 VSS.n666 585
R974 VSS.n2113 VSS.n2112 585
R975 VSS.n2114 VSS.n2113 585
R976 VSS.n664 VSS.n663 585
R977 VSS.n2115 VSS.n664 585
R978 VSS.n2118 VSS.n2117 585
R979 VSS.n2117 VSS.n2116 585
R980 VSS.n2119 VSS.n662 585
R981 VSS.n665 VSS.n662 585
R982 VSS.n2121 VSS.n2120 585
R983 VSS.n2122 VSS.n2121 585
R984 VSS.n312 VSS.n311 585
R985 VSS.n315 VSS.n312 585
R986 VSS.n2133 VSS.n2132 585
R987 VSS.n2132 VSS.n2131 585
R988 VSS.n2134 VSS.n309 585
R989 VSS.n655 VSS.n309 585
R990 VSS.n2136 VSS.n2135 585
R991 VSS.n2137 VSS.n2136 585
R992 VSS.n310 VSS.n308 585
R993 VSS.n308 VSS.n305 585
R994 VSS.n297 VSS.n296 585
R995 VSS.n299 VSS.n297 585
R996 VSS.n2147 VSS.n2146 585
R997 VSS.n2146 VSS.n2145 585
R998 VSS.n2148 VSS.n294 585
R999 VSS.n644 VSS.n294 585
R1000 VSS.n2150 VSS.n2149 585
R1001 VSS.n2151 VSS.n2150 585
R1002 VSS.n295 VSS.n293 585
R1003 VSS.n293 VSS.n290 585
R1004 VSS.n281 VSS.n280 585
R1005 VSS.n637 VSS.n281 585
R1006 VSS.n2161 VSS.n2160 585
R1007 VSS.n2160 VSS.n2159 585
R1008 VSS.n2162 VSS.n278 585
R1009 VSS.n282 VSS.n278 585
R1010 VSS.n2164 VSS.n2163 585
R1011 VSS.n2165 VSS.n2164 585
R1012 VSS.n279 VSS.n277 585
R1013 VSS.n277 VSS.n274 585
R1014 VSS.n264 VSS.n263 585
R1015 VSS.n268 VSS.n264 585
R1016 VSS.n2175 VSS.n2174 585
R1017 VSS.n2174 VSS.n2173 585
R1018 VSS.n2176 VSS.n261 585
R1019 VSS.n265 VSS.n261 585
R1020 VSS.n2178 VSS.n2177 585
R1021 VSS.n2179 VSS.n2178 585
R1022 VSS.n262 VSS.n260 585
R1023 VSS.n260 VSS.n257 585
R1024 VSS.n247 VSS.n246 585
R1025 VSS.n249 VSS.n247 585
R1026 VSS.n2189 VSS.n2188 585
R1027 VSS.n2188 VSS.n2187 585
R1028 VSS.n2190 VSS.n244 585
R1029 VSS.n614 VSS.n244 585
R1030 VSS.n2192 VSS.n2191 585
R1031 VSS.n2193 VSS.n2192 585
R1032 VSS.n245 VSS.n243 585
R1033 VSS.n1966 VSS.n1965 585
R1034 VSS.n1968 VSS.n1967 585
R1035 VSS.n1970 VSS.n1962 585
R1036 VSS.n1972 VSS.n1971 585
R1037 VSS.n1973 VSS.n1904 585
R1038 VSS.n1207 VSS.n1206 585
R1039 VSS.n1208 VSS.n1207 585
R1040 VSS.n820 VSS.n819 585
R1041 VSS.n1209 VSS.n820 585
R1042 VSS.n1219 VSS.n1218 585
R1043 VSS.n1218 VSS.n1217 585
R1044 VSS.n1220 VSS.n818 585
R1045 VSS.n822 VSS.n818 585
R1046 VSS.n1222 VSS.n1221 585
R1047 VSS.n1223 VSS.n1222 585
R1048 VSS.n813 VSS.n812 585
R1049 VSS.n1224 VSS.n813 585
R1050 VSS.n1233 VSS.n1232 585
R1051 VSS.n1232 VSS.n1231 585
R1052 VSS.n1234 VSS.n811 585
R1053 VSS.n811 VSS.n809 585
R1054 VSS.n1236 VSS.n1235 585
R1055 VSS.n1237 VSS.n1236 585
R1056 VSS.n805 VSS.n804 585
R1057 VSS.n810 VSS.n805 585
R1058 VSS.n1245 VSS.n1244 585
R1059 VSS.n1244 VSS.n1243 585
R1060 VSS.n1246 VSS.n803 585
R1061 VSS.n803 VSS.n801 585
R1062 VSS.n1248 VSS.n1247 585
R1063 VSS.n1249 VSS.n1248 585
R1064 VSS.n797 VSS.n796 585
R1065 VSS.n802 VSS.n797 585
R1066 VSS.n1257 VSS.n1256 585
R1067 VSS.n1256 VSS.n1255 585
R1068 VSS.n1258 VSS.n795 585
R1069 VSS.n795 VSS.n793 585
R1070 VSS.n1260 VSS.n1259 585
R1071 VSS.n1261 VSS.n1260 585
R1072 VSS.n789 VSS.n788 585
R1073 VSS.n794 VSS.n789 585
R1074 VSS.n1269 VSS.n1268 585
R1075 VSS.n1268 VSS.n1267 585
R1076 VSS.n1270 VSS.n787 585
R1077 VSS.n787 VSS.n786 585
R1078 VSS.n1272 VSS.n1271 585
R1079 VSS.n1273 VSS.n1272 585
R1080 VSS.n781 VSS.n780 585
R1081 VSS.n782 VSS.n781 585
R1082 VSS.n1281 VSS.n1280 585
R1083 VSS.n1280 VSS.n1279 585
R1084 VSS.n1282 VSS.n779 585
R1085 VSS.n779 VSS.n778 585
R1086 VSS.n1284 VSS.n1283 585
R1087 VSS.n1285 VSS.n1284 585
R1088 VSS.n773 VSS.n772 585
R1089 VSS.n774 VSS.n773 585
R1090 VSS.n1293 VSS.n1292 585
R1091 VSS.n1292 VSS.n1291 585
R1092 VSS.n1294 VSS.n771 585
R1093 VSS.n771 VSS.n770 585
R1094 VSS.n1296 VSS.n1295 585
R1095 VSS.n1297 VSS.n1296 585
R1096 VSS.n765 VSS.n764 585
R1097 VSS.n766 VSS.n765 585
R1098 VSS.n1305 VSS.n1304 585
R1099 VSS.n1304 VSS.n1303 585
R1100 VSS.n1306 VSS.n763 585
R1101 VSS.n763 VSS.n762 585
R1102 VSS.n1308 VSS.n1307 585
R1103 VSS.n1309 VSS.n1308 585
R1104 VSS.n757 VSS.n756 585
R1105 VSS.n758 VSS.n757 585
R1106 VSS.n1317 VSS.n1316 585
R1107 VSS.n1316 VSS.n1315 585
R1108 VSS.n1318 VSS.n755 585
R1109 VSS.n755 VSS.n754 585
R1110 VSS.n1320 VSS.n1319 585
R1111 VSS.n1321 VSS.n1320 585
R1112 VSS.n749 VSS.n748 585
R1113 VSS.n750 VSS.n749 585
R1114 VSS.n1330 VSS.n1329 585
R1115 VSS.n1329 VSS.n1328 585
R1116 VSS.n1331 VSS.n747 585
R1117 VSS.n1327 VSS.n747 585
R1118 VSS.n1333 VSS.n1332 585
R1119 VSS.n1334 VSS.n1333 585
R1120 VSS.n742 VSS.n741 585
R1121 VSS.n743 VSS.n742 585
R1122 VSS.n1343 VSS.n1342 585
R1123 VSS.n1342 VSS.n1341 585
R1124 VSS.n1344 VSS.n740 585
R1125 VSS.n1340 VSS.n740 585
R1126 VSS.n1346 VSS.n1345 585
R1127 VSS.n1347 VSS.n1346 585
R1128 VSS.n735 VSS.n734 585
R1129 VSS.n736 VSS.n735 585
R1130 VSS.n1356 VSS.n1355 585
R1131 VSS.n1355 VSS.n1354 585
R1132 VSS.n1357 VSS.n733 585
R1133 VSS.n1353 VSS.n733 585
R1134 VSS.n1359 VSS.n1358 585
R1135 VSS.n1360 VSS.n1359 585
R1136 VSS.n728 VSS.n727 585
R1137 VSS.n729 VSS.n728 585
R1138 VSS.n1370 VSS.n1369 585
R1139 VSS.n1369 VSS.n1368 585
R1140 VSS.n1371 VSS.n726 585
R1141 VSS.n1367 VSS.n726 585
R1142 VSS.n1373 VSS.n1372 585
R1143 VSS.n1374 VSS.n1373 585
R1144 VSS.n723 VSS.n722 585
R1145 VSS.n722 VSS.n690 585
R1146 VSS.n1494 VSS.n1493 585
R1147 VSS.n1492 VSS.n721 585
R1148 VSS.n1491 VSS.n720 585
R1149 VSS.n1496 VSS.n720 585
R1150 VSS.n1490 VSS.n1489 585
R1151 VSS.n1488 VSS.n1487 585
R1152 VSS.n1486 VSS.n1485 585
R1153 VSS.n1484 VSS.n1483 585
R1154 VSS.n1482 VSS.n1481 585
R1155 VSS.n1480 VSS.n1479 585
R1156 VSS.n1478 VSS.n1477 585
R1157 VSS.n1476 VSS.n1475 585
R1158 VSS.n1474 VSS.n1473 585
R1159 VSS.n1472 VSS.n1471 585
R1160 VSS.n1470 VSS.n1469 585
R1161 VSS.n1468 VSS.n1467 585
R1162 VSS.n1466 VSS.n1465 585
R1163 VSS.n1464 VSS.n1463 585
R1164 VSS.n1462 VSS.n1461 585
R1165 VSS.n1460 VSS.n1459 585
R1166 VSS.n1458 VSS.n1457 585
R1167 VSS.n1456 VSS.n1455 585
R1168 VSS.n1454 VSS.n1453 585
R1169 VSS.n1452 VSS.n1451 585
R1170 VSS.n1450 VSS.n1449 585
R1171 VSS.n1448 VSS.n1447 585
R1172 VSS.n1446 VSS.n1445 585
R1173 VSS.n1444 VSS.n1443 585
R1174 VSS.n1442 VSS.n1441 585
R1175 VSS.n1440 VSS.n1439 585
R1176 VSS.n1438 VSS.n1437 585
R1177 VSS.n1436 VSS.n1435 585
R1178 VSS.n1434 VSS.n1433 585
R1179 VSS.n1432 VSS.n1431 585
R1180 VSS.n1430 VSS.n1429 585
R1181 VSS.n1428 VSS.n1427 585
R1182 VSS.n1426 VSS.n1425 585
R1183 VSS.n1424 VSS.n1423 585
R1184 VSS.n1422 VSS.n1421 585
R1185 VSS.n1420 VSS.n1419 585
R1186 VSS.n1418 VSS.n1417 585
R1187 VSS.n1416 VSS.n1415 585
R1188 VSS.n1414 VSS.n1413 585
R1189 VSS.n1412 VSS.n1411 585
R1190 VSS.n1410 VSS.n1409 585
R1191 VSS.n1408 VSS.n1407 585
R1192 VSS.n1406 VSS.n1405 585
R1193 VSS.n1404 VSS.n1403 585
R1194 VSS.n1402 VSS.n1401 585
R1195 VSS.n1400 VSS.n1399 585
R1196 VSS.n1398 VSS.n1397 585
R1197 VSS.n1396 VSS.n1395 585
R1198 VSS.n1394 VSS.n1393 585
R1199 VSS.n1392 VSS.n1391 585
R1200 VSS.n1390 VSS.n1389 585
R1201 VSS.n1388 VSS.n1387 585
R1202 VSS.n1386 VSS.n1385 585
R1203 VSS.n1384 VSS.n1383 585
R1204 VSS.n1382 VSS.n1381 585
R1205 VSS.n1380 VSS.n1379 585
R1206 VSS.n1378 VSS.n719 585
R1207 VSS.n1496 VSS.n719 585
R1208 VSS.n1377 VSS.n1376 585
R1209 VSS.n1376 VSS.n690 585
R1210 VSS.n1375 VSS.n724 585
R1211 VSS.n1375 VSS.n1374 585
R1212 VSS.n1364 VSS.n725 585
R1213 VSS.n1367 VSS.n725 585
R1214 VSS.n1366 VSS.n1365 585
R1215 VSS.n1368 VSS.n1366 585
R1216 VSS.n1363 VSS.n730 585
R1217 VSS.n730 VSS.n729 585
R1218 VSS.n1362 VSS.n1361 585
R1219 VSS.n1361 VSS.n1360 585
R1220 VSS.n732 VSS.n731 585
R1221 VSS.n1353 VSS.n732 585
R1222 VSS.n1352 VSS.n1351 585
R1223 VSS.n1354 VSS.n1352 585
R1224 VSS.n1350 VSS.n737 585
R1225 VSS.n737 VSS.n736 585
R1226 VSS.n1349 VSS.n1348 585
R1227 VSS.n1348 VSS.n1347 585
R1228 VSS.n739 VSS.n738 585
R1229 VSS.n1340 VSS.n739 585
R1230 VSS.n1339 VSS.n1338 585
R1231 VSS.n1341 VSS.n1339 585
R1232 VSS.n1337 VSS.n744 585
R1233 VSS.n744 VSS.n743 585
R1234 VSS.n1336 VSS.n1335 585
R1235 VSS.n1335 VSS.n1334 585
R1236 VSS.n746 VSS.n745 585
R1237 VSS.n1327 VSS.n746 585
R1238 VSS.n1326 VSS.n1325 585
R1239 VSS.n1328 VSS.n1326 585
R1240 VSS.n1324 VSS.n751 585
R1241 VSS.n751 VSS.n750 585
R1242 VSS.n1323 VSS.n1322 585
R1243 VSS.n1322 VSS.n1321 585
R1244 VSS.n753 VSS.n752 585
R1245 VSS.n754 VSS.n753 585
R1246 VSS.n1314 VSS.n1313 585
R1247 VSS.n1315 VSS.n1314 585
R1248 VSS.n1312 VSS.n759 585
R1249 VSS.n759 VSS.n758 585
R1250 VSS.n1311 VSS.n1310 585
R1251 VSS.n1310 VSS.n1309 585
R1252 VSS.n761 VSS.n760 585
R1253 VSS.n762 VSS.n761 585
R1254 VSS.n1302 VSS.n1301 585
R1255 VSS.n1303 VSS.n1302 585
R1256 VSS.n1300 VSS.n767 585
R1257 VSS.n767 VSS.n766 585
R1258 VSS.n1299 VSS.n1298 585
R1259 VSS.n1298 VSS.n1297 585
R1260 VSS.n769 VSS.n768 585
R1261 VSS.n770 VSS.n769 585
R1262 VSS.n1290 VSS.n1289 585
R1263 VSS.n1291 VSS.n1290 585
R1264 VSS.n1288 VSS.n775 585
R1265 VSS.n775 VSS.n774 585
R1266 VSS.n1287 VSS.n1286 585
R1267 VSS.n1286 VSS.n1285 585
R1268 VSS.n777 VSS.n776 585
R1269 VSS.n778 VSS.n777 585
R1270 VSS.n1278 VSS.n1277 585
R1271 VSS.n1279 VSS.n1278 585
R1272 VSS.n1276 VSS.n783 585
R1273 VSS.n783 VSS.n782 585
R1274 VSS.n1275 VSS.n1274 585
R1275 VSS.n1274 VSS.n1273 585
R1276 VSS.n785 VSS.n784 585
R1277 VSS.n786 VSS.n785 585
R1278 VSS.n1266 VSS.n1265 585
R1279 VSS.n1267 VSS.n1266 585
R1280 VSS.n1264 VSS.n790 585
R1281 VSS.n794 VSS.n790 585
R1282 VSS.n1263 VSS.n1262 585
R1283 VSS.n1262 VSS.n1261 585
R1284 VSS.n792 VSS.n791 585
R1285 VSS.n793 VSS.n792 585
R1286 VSS.n1254 VSS.n1253 585
R1287 VSS.n1255 VSS.n1254 585
R1288 VSS.n1252 VSS.n798 585
R1289 VSS.n802 VSS.n798 585
R1290 VSS.n1251 VSS.n1250 585
R1291 VSS.n1250 VSS.n1249 585
R1292 VSS.n800 VSS.n799 585
R1293 VSS.n801 VSS.n800 585
R1294 VSS.n1242 VSS.n1241 585
R1295 VSS.n1243 VSS.n1242 585
R1296 VSS.n1240 VSS.n806 585
R1297 VSS.n810 VSS.n806 585
R1298 VSS.n1239 VSS.n1238 585
R1299 VSS.n1238 VSS.n1237 585
R1300 VSS.n808 VSS.n807 585
R1301 VSS.n809 VSS.n808 585
R1302 VSS.n1230 VSS.n1229 585
R1303 VSS.n1231 VSS.n1230 585
R1304 VSS.n1228 VSS.n814 585
R1305 VSS.n1224 VSS.n814 585
R1306 VSS.n1227 VSS.n1226 585
R1307 VSS.n1226 VSS.n1225 585
R1308 VSS.n816 VSS.n815 585
R1309 VSS.n817 VSS.n816 585
R1310 VSS.n1215 VSS.n1214 585
R1311 VSS.n1216 VSS.n1215 585
R1312 VSS.n1213 VSS.n823 585
R1313 VSS.n823 VSS.n821 585
R1314 VSS.n1212 VSS.n1211 585
R1315 VSS.n1211 VSS.n1210 585
R1316 VSS.n825 VSS.n824 585
R1317 VSS.n1104 VSS.n1101 585
R1318 VSS.n1106 VSS.n1105 585
R1319 VSS.n1107 VSS.n868 585
R1320 VSS.n1109 VSS.n1108 585
R1321 VSS.n1111 VSS.n866 585
R1322 VSS.n1113 VSS.n1112 585
R1323 VSS.n1114 VSS.n865 585
R1324 VSS.n1116 VSS.n1115 585
R1325 VSS.n1118 VSS.n863 585
R1326 VSS.n1120 VSS.n1119 585
R1327 VSS.n1121 VSS.n862 585
R1328 VSS.n1123 VSS.n1122 585
R1329 VSS.n1125 VSS.n860 585
R1330 VSS.n1127 VSS.n1126 585
R1331 VSS.n1128 VSS.n859 585
R1332 VSS.n1130 VSS.n1129 585
R1333 VSS.n1132 VSS.n857 585
R1334 VSS.n1134 VSS.n1133 585
R1335 VSS.n1135 VSS.n856 585
R1336 VSS.n1137 VSS.n1136 585
R1337 VSS.n1139 VSS.n854 585
R1338 VSS.n1141 VSS.n1140 585
R1339 VSS.n1142 VSS.n853 585
R1340 VSS.n1144 VSS.n1143 585
R1341 VSS.n1146 VSS.n851 585
R1342 VSS.n1148 VSS.n1147 585
R1343 VSS.n1149 VSS.n850 585
R1344 VSS.n1151 VSS.n1150 585
R1345 VSS.n1153 VSS.n848 585
R1346 VSS.n1155 VSS.n1154 585
R1347 VSS.n1156 VSS.n847 585
R1348 VSS.n1158 VSS.n1157 585
R1349 VSS.n1160 VSS.n845 585
R1350 VSS.n1162 VSS.n1161 585
R1351 VSS.n1163 VSS.n844 585
R1352 VSS.n1165 VSS.n1164 585
R1353 VSS.n1167 VSS.n842 585
R1354 VSS.n1169 VSS.n1168 585
R1355 VSS.n1170 VSS.n841 585
R1356 VSS.n1172 VSS.n1171 585
R1357 VSS.n1174 VSS.n839 585
R1358 VSS.n1176 VSS.n1175 585
R1359 VSS.n1177 VSS.n838 585
R1360 VSS.n1179 VSS.n1178 585
R1361 VSS.n1181 VSS.n836 585
R1362 VSS.n1183 VSS.n1182 585
R1363 VSS.n1184 VSS.n835 585
R1364 VSS.n1186 VSS.n1185 585
R1365 VSS.n1188 VSS.n833 585
R1366 VSS.n1190 VSS.n1189 585
R1367 VSS.n1191 VSS.n832 585
R1368 VSS.n1193 VSS.n1192 585
R1369 VSS.n1195 VSS.n830 585
R1370 VSS.n1197 VSS.n1196 585
R1371 VSS.n1198 VSS.n829 585
R1372 VSS.n1200 VSS.n1199 585
R1373 VSS.n1202 VSS.n827 585
R1374 VSS.n1204 VSS.n1203 585
R1375 VSS.n1205 VSS.n826 585
R1376 VSS.n1787 VSS.n1617 533.088
R1377 VSS.n1775 VSS.n1615 533.088
R1378 VSS.n2107 VSS.n671 504.736
R1379 VSS.n1222 VSS.n813 463.529
R1380 VSS.n2224 VSS.n214 394
R1381 VSS.n2220 VSS.n214 394
R1382 VSS.n2220 VSS.n217 394
R1383 VSS.n2216 VSS.n217 394
R1384 VSS.n2216 VSS.n222 394
R1385 VSS.n2212 VSS.n222 394
R1386 VSS.n2212 VSS.n224 394
R1387 VSS.n2208 VSS.n224 394
R1388 VSS.n2208 VSS.n229 394
R1389 VSS.n2204 VSS.n229 394
R1390 VSS.n2204 VSS.n231 394
R1391 VSS.n2200 VSS.n231 394
R1392 VSS.n2200 VSS.n236 394
R1393 VSS.n2196 VSS.n236 394
R1394 VSS.n2196 VSS.n238 394
R1395 VSS.n252 VSS.n238 394
R1396 VSS.n252 VSS.n250 394
R1397 VSS.n2185 VSS.n250 394
R1398 VSS.n2185 VSS.n251 394
R1399 VSS.n2181 VSS.n251 394
R1400 VSS.n2181 VSS.n256 394
R1401 VSS.n269 VSS.n256 394
R1402 VSS.n2171 VSS.n269 394
R1403 VSS.n2171 VSS.n270 394
R1404 VSS.n2167 VSS.n270 394
R1405 VSS.n2167 VSS.n273 394
R1406 VSS.n285 VSS.n273 394
R1407 VSS.n2157 VSS.n285 394
R1408 VSS.n2157 VSS.n286 394
R1409 VSS.n2153 VSS.n286 394
R1410 VSS.n2153 VSS.n289 394
R1411 VSS.n300 VSS.n289 394
R1412 VSS.n2143 VSS.n300 394
R1413 VSS.n2143 VSS.n301 394
R1414 VSS.n2139 VSS.n301 394
R1415 VSS.n2139 VSS.n304 394
R1416 VSS.n316 VSS.n304 394
R1417 VSS.n2129 VSS.n316 394
R1418 VSS.n504 VSS.n503 394
R1419 VSS.n508 VSS.n507 394
R1420 VSS.n512 VSS.n511 394
R1421 VSS.n516 VSS.n515 394
R1422 VSS.n520 VSS.n519 394
R1423 VSS.n528 VSS.n527 394
R1424 VSS.n532 VSS.n531 394
R1425 VSS.n536 VSS.n535 394
R1426 VSS.n540 VSS.n539 394
R1427 VSS.n544 VSS.n543 394
R1428 VSS.n548 VSS.n547 394
R1429 VSS.n552 VSS.n551 394
R1430 VSS.n556 VSS.n555 394
R1431 VSS.n560 VSS.n559 394
R1432 VSS.n564 VSS.n563 394
R1433 VSS.n572 VSS.n571 394
R1434 VSS.n576 VSS.n575 394
R1435 VSS.n580 VSS.n579 394
R1436 VSS.n584 VSS.n583 394
R1437 VSS.n588 VSS.n587 394
R1438 VSS.n593 VSS.n211 394
R1439 VSS.n593 VSS.n218 394
R1440 VSS.n219 VSS.n218 394
R1441 VSS.n220 VSS.n219 394
R1442 VSS.n598 VSS.n220 394
R1443 VSS.n598 VSS.n225 394
R1444 VSS.n226 VSS.n225 394
R1445 VSS.n227 VSS.n226 394
R1446 VSS.n603 VSS.n227 394
R1447 VSS.n603 VSS.n232 394
R1448 VSS.n233 VSS.n232 394
R1449 VSS.n234 VSS.n233 394
R1450 VSS.n608 VSS.n234 394
R1451 VSS.n608 VSS.n240 394
R1452 VSS.n241 VSS.n240 394
R1453 VSS.n613 VSS.n241 394
R1454 VSS.n616 VSS.n613 394
R1455 VSS.n616 VSS.n248 394
R1456 VSS.n620 VSS.n248 394
R1457 VSS.n620 VSS.n258 394
R1458 VSS.n624 VSS.n258 394
R1459 VSS.n625 VSS.n624 394
R1460 VSS.n625 VSS.n267 394
R1461 VSS.n629 VSS.n267 394
R1462 VSS.n629 VSS.n275 394
R1463 VSS.n633 VSS.n275 394
R1464 VSS.n634 VSS.n633 394
R1465 VSS.n634 VSS.n284 394
R1466 VSS.n639 VSS.n284 394
R1467 VSS.n639 VSS.n291 394
R1468 VSS.n643 VSS.n291 394
R1469 VSS.n646 VSS.n643 394
R1470 VSS.n646 VSS.n298 394
R1471 VSS.n650 VSS.n298 394
R1472 VSS.n650 VSS.n306 394
R1473 VSS.n654 VSS.n306 394
R1474 VSS.n657 VSS.n654 394
R1475 VSS.n657 VSS.n314 394
R1476 VSS.n2125 VSS.n320 394
R1477 VSS.n344 VSS.n320 394
R1478 VSS.n348 VSS.n347 394
R1479 VSS.n352 VSS.n351 394
R1480 VSS.n356 VSS.n355 394
R1481 VSS.n360 VSS.n359 394
R1482 VSS.n364 VSS.n363 394
R1483 VSS.n368 VSS.n367 394
R1484 VSS.n372 VSS.n371 394
R1485 VSS.n376 VSS.n375 394
R1486 VSS.n380 VSS.n379 394
R1487 VSS.n384 VSS.n383 394
R1488 VSS.n388 VSS.n387 394
R1489 VSS.n392 VSS.n391 394
R1490 VSS.n396 VSS.n395 394
R1491 VSS.n400 VSS.n399 394
R1492 VSS.n404 VSS.n403 394
R1493 VSS.n408 VSS.n407 394
R1494 VSS.n412 VSS.n411 394
R1495 VSS.n416 VSS.n415 394
R1496 VSS.n420 VSS.n419 394
R1497 VSS.n424 VSS.n423 394
R1498 VSS.n428 VSS.n427 394
R1499 VSS.n661 VSS.n343 394
R1500 VSS.n1980 VSS.n1529 394
R1501 VSS.n1980 VSS.n1527 394
R1502 VSS.n1984 VSS.n1527 394
R1503 VSS.n1984 VSS.n1525 394
R1504 VSS.n1988 VSS.n1525 394
R1505 VSS.n1988 VSS.n1523 394
R1506 VSS.n1992 VSS.n1523 394
R1507 VSS.n1992 VSS.n1521 394
R1508 VSS.n1996 VSS.n1521 394
R1509 VSS.n1996 VSS.n1519 394
R1510 VSS.n2000 VSS.n1519 394
R1511 VSS.n2000 VSS.n1517 394
R1512 VSS.n2004 VSS.n1517 394
R1513 VSS.n2004 VSS.n1515 394
R1514 VSS.n2008 VSS.n1515 394
R1515 VSS.n2008 VSS.n1513 394
R1516 VSS.n2012 VSS.n1513 394
R1517 VSS.n2012 VSS.n1511 394
R1518 VSS.n2016 VSS.n1511 394
R1519 VSS.n2016 VSS.n1509 394
R1520 VSS.n2020 VSS.n1509 394
R1521 VSS.n2020 VSS.n1507 394
R1522 VSS.n2024 VSS.n1507 394
R1523 VSS.n2024 VSS.n1505 394
R1524 VSS.n2028 VSS.n1505 394
R1525 VSS.n2028 VSS.n1503 394
R1526 VSS.n2032 VSS.n1503 394
R1527 VSS.n2032 VSS.n1501 394
R1528 VSS.n2036 VSS.n1501 394
R1529 VSS.n2036 VSS.n1499 394
R1530 VSS.n1909 VSS.n1908 394
R1531 VSS.n1913 VSS.n1912 394
R1532 VSS.n1917 VSS.n1916 394
R1533 VSS.n1921 VSS.n1920 394
R1534 VSS.n1925 VSS.n1924 394
R1535 VSS.n1929 VSS.n1928 394
R1536 VSS.n1933 VSS.n1932 394
R1537 VSS.n1937 VSS.n1936 394
R1538 VSS.n1941 VSS.n1940 394
R1539 VSS.n1945 VSS.n1944 394
R1540 VSS.n1949 VSS.n1948 394
R1541 VSS.n1953 VSS.n1952 394
R1542 VSS.n1957 VSS.n1956 394
R1543 VSS.n1959 VSS.n1903 394
R1544 VSS.n1975 VSS.n1904 394
R1545 VSS.n1971 VSS.n1970 394
R1546 VSS.n1968 VSS.n1965 394
R1547 VSS.n2192 VSS.n244 394
R1548 VSS.n2188 VSS.n244 394
R1549 VSS.n2188 VSS.n247 394
R1550 VSS.n260 VSS.n247 394
R1551 VSS.n2178 VSS.n260 394
R1552 VSS.n2178 VSS.n261 394
R1553 VSS.n2174 VSS.n261 394
R1554 VSS.n2174 VSS.n264 394
R1555 VSS.n277 VSS.n264 394
R1556 VSS.n2164 VSS.n277 394
R1557 VSS.n2164 VSS.n278 394
R1558 VSS.n2160 VSS.n278 394
R1559 VSS.n2160 VSS.n281 394
R1560 VSS.n293 VSS.n281 394
R1561 VSS.n2150 VSS.n293 394
R1562 VSS.n2150 VSS.n294 394
R1563 VSS.n2146 VSS.n294 394
R1564 VSS.n2146 VSS.n297 394
R1565 VSS.n308 VSS.n297 394
R1566 VSS.n2136 VSS.n308 394
R1567 VSS.n2136 VSS.n309 394
R1568 VSS.n2132 VSS.n309 394
R1569 VSS.n2132 VSS.n312 394
R1570 VSS.n2121 VSS.n312 394
R1571 VSS.n2121 VSS.n662 394
R1572 VSS.n2117 VSS.n662 394
R1573 VSS.n2117 VSS.n664 394
R1574 VSS.n2113 VSS.n664 394
R1575 VSS.n2113 VSS.n666 394
R1576 VSS.n2109 VSS.n666 394
R1577 VSS.n1498 VSS.n1497 394
R1578 VSS.n2085 VSS.n1497 394
R1579 VSS.n2083 VSS.n2082 394
R1580 VSS.n2079 VSS.n2078 394
R1581 VSS.n2075 VSS.n2074 394
R1582 VSS.n2071 VSS.n2070 394
R1583 VSS.n2067 VSS.n2066 394
R1584 VSS.n2063 VSS.n2062 394
R1585 VSS.n2059 VSS.n2058 394
R1586 VSS.n2055 VSS.n2054 394
R1587 VSS.n2051 VSS.n2050 394
R1588 VSS.n2047 VSS.n2046 394
R1589 VSS.n2043 VSS.n2042 394
R1590 VSS.n2039 VSS.n676 394
R1591 VSS.n2094 VSS.n674 394
R1592 VSS.n2105 VSS.n674 394
R1593 VSS.n673 VSS.n672 394
R1594 VSS.n2100 VSS.n672 394
R1595 VSS.n2098 VSS.n668 394
R1596 VSS.n1875 VSS.n1534 394
R1597 VSS.n1875 VSS.n1540 394
R1598 VSS.n1871 VSS.n1540 394
R1599 VSS.n1871 VSS.n1542 394
R1600 VSS.n1867 VSS.n1542 394
R1601 VSS.n1867 VSS.n1547 394
R1602 VSS.n1863 VSS.n1547 394
R1603 VSS.n1863 VSS.n1549 394
R1604 VSS.n1859 VSS.n1549 394
R1605 VSS.n1859 VSS.n1554 394
R1606 VSS.n1855 VSS.n1554 394
R1607 VSS.n1855 VSS.n1556 394
R1608 VSS.n1851 VSS.n1556 394
R1609 VSS.n1851 VSS.n1561 394
R1610 VSS.n1847 VSS.n1561 394
R1611 VSS.n1847 VSS.n1563 394
R1612 VSS.n1843 VSS.n1563 394
R1613 VSS.n1843 VSS.n1568 394
R1614 VSS.n1839 VSS.n1568 394
R1615 VSS.n1839 VSS.n1570 394
R1616 VSS.n1835 VSS.n1570 394
R1617 VSS.n1835 VSS.n1575 394
R1618 VSS.n1831 VSS.n1575 394
R1619 VSS.n1831 VSS.n1577 394
R1620 VSS.n1827 VSS.n1577 394
R1621 VSS.n1827 VSS.n1582 394
R1622 VSS.n1823 VSS.n1582 394
R1623 VSS.n1823 VSS.n1584 394
R1624 VSS.n1819 VSS.n1584 394
R1625 VSS.n1819 VSS.n1589 394
R1626 VSS.n1815 VSS.n1589 394
R1627 VSS.n1815 VSS.n1591 394
R1628 VSS.n1811 VSS.n1591 394
R1629 VSS.n1811 VSS.n1596 394
R1630 VSS.n1807 VSS.n1596 394
R1631 VSS.n1807 VSS.n1598 394
R1632 VSS.n1803 VSS.n1598 394
R1633 VSS.n1803 VSS.n1603 394
R1634 VSS.n1799 VSS.n1603 394
R1635 VSS.n1799 VSS.n1605 394
R1636 VSS.n1795 VSS.n1605 394
R1637 VSS.n1795 VSS.n1610 394
R1638 VSS.n1791 VSS.n1610 394
R1639 VSS.n1791 VSS.n1612 394
R1640 VSS.n1787 VSS.n1612 394
R1641 VSS.n1533 VSS.n1532 394
R1642 VSS.n1881 VSS.n1532 394
R1643 VSS.n1878 VSS.n1877 394
R1644 VSS.n1877 VSS.n1537 394
R1645 VSS.n1543 VSS.n1537 394
R1646 VSS.n1544 VSS.n1543 394
R1647 VSS.n1545 VSS.n1544 394
R1648 VSS.n1725 VSS.n1545 394
R1649 VSS.n1725 VSS.n1550 394
R1650 VSS.n1551 VSS.n1550 394
R1651 VSS.n1552 VSS.n1551 394
R1652 VSS.n1730 VSS.n1552 394
R1653 VSS.n1730 VSS.n1557 394
R1654 VSS.n1558 VSS.n1557 394
R1655 VSS.n1559 VSS.n1558 394
R1656 VSS.n1735 VSS.n1559 394
R1657 VSS.n1735 VSS.n1564 394
R1658 VSS.n1565 VSS.n1564 394
R1659 VSS.n1566 VSS.n1565 394
R1660 VSS.n1740 VSS.n1566 394
R1661 VSS.n1740 VSS.n1571 394
R1662 VSS.n1572 VSS.n1571 394
R1663 VSS.n1573 VSS.n1572 394
R1664 VSS.n1745 VSS.n1573 394
R1665 VSS.n1745 VSS.n1578 394
R1666 VSS.n1579 VSS.n1578 394
R1667 VSS.n1580 VSS.n1579 394
R1668 VSS.n1750 VSS.n1580 394
R1669 VSS.n1750 VSS.n1585 394
R1670 VSS.n1586 VSS.n1585 394
R1671 VSS.n1587 VSS.n1586 394
R1672 VSS.n1755 VSS.n1587 394
R1673 VSS.n1755 VSS.n1592 394
R1674 VSS.n1593 VSS.n1592 394
R1675 VSS.n1594 VSS.n1593 394
R1676 VSS.n1760 VSS.n1594 394
R1677 VSS.n1760 VSS.n1599 394
R1678 VSS.n1600 VSS.n1599 394
R1679 VSS.n1601 VSS.n1600 394
R1680 VSS.n1765 VSS.n1601 394
R1681 VSS.n1765 VSS.n1606 394
R1682 VSS.n1607 VSS.n1606 394
R1683 VSS.n1608 VSS.n1607 394
R1684 VSS.n1770 VSS.n1608 394
R1685 VSS.n1770 VSS.n1613 394
R1686 VSS.n1614 VSS.n1613 394
R1687 VSS.n1615 VSS.n1614 394
R1688 VSS.n2381 VSS.n127 394
R1689 VSS.n2381 VSS.n128 394
R1690 VSS.n2377 VSS.n128 394
R1691 VSS.n2377 VSS.n131 394
R1692 VSS.n2373 VSS.n131 394
R1693 VSS.n2373 VSS.n136 394
R1694 VSS.n2369 VSS.n136 394
R1695 VSS.n2369 VSS.n138 394
R1696 VSS.n2365 VSS.n138 394
R1697 VSS.n2365 VSS.n142 394
R1698 VSS.n2361 VSS.n142 394
R1699 VSS.n2361 VSS.n144 394
R1700 VSS.n2357 VSS.n144 394
R1701 VSS.n2357 VSS.n149 394
R1702 VSS.n2353 VSS.n149 394
R1703 VSS.n2353 VSS.n151 394
R1704 VSS.n2349 VSS.n151 394
R1705 VSS.n2349 VSS.n156 394
R1706 VSS.n2345 VSS.n156 394
R1707 VSS.n2345 VSS.n158 394
R1708 VSS.n2341 VSS.n158 394
R1709 VSS.n2341 VSS.n163 394
R1710 VSS.n2337 VSS.n163 394
R1711 VSS.n1643 VSS.n1642 394
R1712 VSS.n1647 VSS.n1646 394
R1713 VSS.n1651 VSS.n1650 394
R1714 VSS.n1655 VSS.n1654 394
R1715 VSS.n1659 VSS.n1658 394
R1716 VSS.n1667 VSS.n1666 394
R1717 VSS.n1671 VSS.n1670 394
R1718 VSS.n1675 VSS.n1674 394
R1719 VSS.n1679 VSS.n1678 394
R1720 VSS.n1683 VSS.n1682 394
R1721 VSS.n1687 VSS.n1686 394
R1722 VSS.n1691 VSS.n1690 394
R1723 VSS.n1695 VSS.n1694 394
R1724 VSS.n1699 VSS.n1698 394
R1725 VSS.n1703 VSS.n1702 394
R1726 VSS.n1711 VSS.n1710 394
R1727 VSS.n1715 VSS.n1638 394
R1728 VSS.n2383 VSS.n124 394
R1729 VSS.n132 VSS.n124 394
R1730 VSS.n133 VSS.n132 394
R1731 VSS.n134 VSS.n133 394
R1732 VSS.n2231 VSS.n134 394
R1733 VSS.n2231 VSS.n139 394
R1734 VSS.n140 VSS.n139 394
R1735 VSS.n141 VSS.n140 394
R1736 VSS.n2236 VSS.n141 394
R1737 VSS.n2236 VSS.n146 394
R1738 VSS.n147 VSS.n146 394
R1739 VSS.n148 VSS.n147 394
R1740 VSS.n2241 VSS.n148 394
R1741 VSS.n2241 VSS.n153 394
R1742 VSS.n154 VSS.n153 394
R1743 VSS.n155 VSS.n154 394
R1744 VSS.n2246 VSS.n155 394
R1745 VSS.n2246 VSS.n160 394
R1746 VSS.n161 VSS.n160 394
R1747 VSS.n162 VSS.n161 394
R1748 VSS.n2251 VSS.n162 394
R1749 VSS.n2251 VSS.n167 394
R1750 VSS.n2333 VSS.n2227 394
R1751 VSS.n2329 VSS.n2227 394
R1752 VSS.n2327 VSS.n2326 394
R1753 VSS.n2323 VSS.n2322 394
R1754 VSS.n2319 VSS.n2318 394
R1755 VSS.n2315 VSS.n2314 394
R1756 VSS.n2311 VSS.n2310 394
R1757 VSS.n2307 VSS.n2306 394
R1758 VSS.n2303 VSS.n2302 394
R1759 VSS.n2299 VSS.n2298 394
R1760 VSS.n2295 VSS.n2294 394
R1761 VSS.n2291 VSS.n2290 394
R1762 VSS.n2287 VSS.n2286 394
R1763 VSS.n2283 VSS.n2282 394
R1764 VSS.n2279 VSS.n2278 394
R1765 VSS.n2275 VSS.n2274 394
R1766 VSS.n2271 VSS.n2270 394
R1767 VSS.n2267 VSS.n2266 394
R1768 VSS.n2263 VSS.n2262 394
R1769 VSS.n2259 VSS.n2258 394
R1770 VSS.n2255 VSS.n187 394
R1771 VSS.n721 VSS.n720 394
R1772 VSS.n1489 VSS.n720 394
R1773 VSS.n1487 VSS.n1486 394
R1774 VSS.n1483 VSS.n1482 394
R1775 VSS.n1479 VSS.n1478 394
R1776 VSS.n1475 VSS.n1474 394
R1777 VSS.n1471 VSS.n1470 394
R1778 VSS.n1467 VSS.n1466 394
R1779 VSS.n1463 VSS.n1462 394
R1780 VSS.n1459 VSS.n1458 394
R1781 VSS.n1455 VSS.n1454 394
R1782 VSS.n1451 VSS.n1450 394
R1783 VSS.n1447 VSS.n1446 394
R1784 VSS.n1443 VSS.n1442 394
R1785 VSS.n1439 VSS.n1438 394
R1786 VSS.n1435 VSS.n1434 394
R1787 VSS.n1431 VSS.n1430 394
R1788 VSS.n1427 VSS.n1426 394
R1789 VSS.n1423 VSS.n1422 394
R1790 VSS.n1419 VSS.n1418 394
R1791 VSS.n1415 VSS.n1414 394
R1792 VSS.n1411 VSS.n1410 394
R1793 VSS.n1407 VSS.n1406 394
R1794 VSS.n1403 VSS.n1402 394
R1795 VSS.n1399 VSS.n1398 394
R1796 VSS.n1395 VSS.n1394 394
R1797 VSS.n1391 VSS.n1390 394
R1798 VSS.n1387 VSS.n1386 394
R1799 VSS.n1383 VSS.n1382 394
R1800 VSS.n1379 VSS.n719 394
R1801 VSS.n1211 VSS.n823 394
R1802 VSS.n1215 VSS.n823 394
R1803 VSS.n1215 VSS.n816 394
R1804 VSS.n1226 VSS.n816 394
R1805 VSS.n1226 VSS.n814 394
R1806 VSS.n1230 VSS.n814 394
R1807 VSS.n1230 VSS.n808 394
R1808 VSS.n1238 VSS.n808 394
R1809 VSS.n1238 VSS.n806 394
R1810 VSS.n1242 VSS.n806 394
R1811 VSS.n1242 VSS.n800 394
R1812 VSS.n1250 VSS.n800 394
R1813 VSS.n1250 VSS.n798 394
R1814 VSS.n1254 VSS.n798 394
R1815 VSS.n1254 VSS.n792 394
R1816 VSS.n1262 VSS.n792 394
R1817 VSS.n1262 VSS.n790 394
R1818 VSS.n1266 VSS.n790 394
R1819 VSS.n1266 VSS.n785 394
R1820 VSS.n1274 VSS.n785 394
R1821 VSS.n1274 VSS.n783 394
R1822 VSS.n1278 VSS.n783 394
R1823 VSS.n1278 VSS.n777 394
R1824 VSS.n1286 VSS.n777 394
R1825 VSS.n1286 VSS.n775 394
R1826 VSS.n1290 VSS.n775 394
R1827 VSS.n1290 VSS.n769 394
R1828 VSS.n1298 VSS.n769 394
R1829 VSS.n1298 VSS.n767 394
R1830 VSS.n1302 VSS.n767 394
R1831 VSS.n1302 VSS.n761 394
R1832 VSS.n1310 VSS.n761 394
R1833 VSS.n1310 VSS.n759 394
R1834 VSS.n1314 VSS.n759 394
R1835 VSS.n1314 VSS.n753 394
R1836 VSS.n1322 VSS.n753 394
R1837 VSS.n1322 VSS.n751 394
R1838 VSS.n1326 VSS.n751 394
R1839 VSS.n1326 VSS.n746 394
R1840 VSS.n1335 VSS.n746 394
R1841 VSS.n1335 VSS.n744 394
R1842 VSS.n1339 VSS.n744 394
R1843 VSS.n1339 VSS.n739 394
R1844 VSS.n1348 VSS.n739 394
R1845 VSS.n1348 VSS.n737 394
R1846 VSS.n1352 VSS.n737 394
R1847 VSS.n1352 VSS.n732 394
R1848 VSS.n1361 VSS.n732 394
R1849 VSS.n1361 VSS.n730 394
R1850 VSS.n1366 VSS.n730 394
R1851 VSS.n1366 VSS.n725 394
R1852 VSS.n1375 VSS.n725 394
R1853 VSS.n1376 VSS.n1375 394
R1854 VSS.n1203 VSS.n1202 394
R1855 VSS.n1200 VSS.n829 394
R1856 VSS.n1196 VSS.n1195 394
R1857 VSS.n1193 VSS.n832 394
R1858 VSS.n1189 VSS.n1188 394
R1859 VSS.n1186 VSS.n835 394
R1860 VSS.n1182 VSS.n1181 394
R1861 VSS.n1179 VSS.n838 394
R1862 VSS.n1175 VSS.n1174 394
R1863 VSS.n1172 VSS.n841 394
R1864 VSS.n1168 VSS.n1167 394
R1865 VSS.n1165 VSS.n844 394
R1866 VSS.n1161 VSS.n1160 394
R1867 VSS.n1158 VSS.n847 394
R1868 VSS.n1154 VSS.n1153 394
R1869 VSS.n1151 VSS.n850 394
R1870 VSS.n1147 VSS.n1146 394
R1871 VSS.n1144 VSS.n853 394
R1872 VSS.n1140 VSS.n1139 394
R1873 VSS.n1137 VSS.n856 394
R1874 VSS.n1133 VSS.n1132 394
R1875 VSS.n1130 VSS.n859 394
R1876 VSS.n1126 VSS.n1125 394
R1877 VSS.n1123 VSS.n862 394
R1878 VSS.n1119 VSS.n1118 394
R1879 VSS.n1116 VSS.n865 394
R1880 VSS.n1112 VSS.n1111 394
R1881 VSS.n1109 VSS.n868 394
R1882 VSS.n1105 VSS.n1104 394
R1883 VSS.n1207 VSS.n820 394
R1884 VSS.n1218 VSS.n820 394
R1885 VSS.n1218 VSS.n818 394
R1886 VSS.n1222 VSS.n818 394
R1887 VSS.n1232 VSS.n813 394
R1888 VSS.n1232 VSS.n811 394
R1889 VSS.n1236 VSS.n811 394
R1890 VSS.n1236 VSS.n805 394
R1891 VSS.n1244 VSS.n805 394
R1892 VSS.n1244 VSS.n803 394
R1893 VSS.n1248 VSS.n803 394
R1894 VSS.n1248 VSS.n797 394
R1895 VSS.n1256 VSS.n797 394
R1896 VSS.n1256 VSS.n795 394
R1897 VSS.n1260 VSS.n795 394
R1898 VSS.n1260 VSS.n789 394
R1899 VSS.n1268 VSS.n789 394
R1900 VSS.n1268 VSS.n787 394
R1901 VSS.n1272 VSS.n787 394
R1902 VSS.n1272 VSS.n781 394
R1903 VSS.n1280 VSS.n781 394
R1904 VSS.n1280 VSS.n779 394
R1905 VSS.n1284 VSS.n779 394
R1906 VSS.n1284 VSS.n773 394
R1907 VSS.n1292 VSS.n773 394
R1908 VSS.n1292 VSS.n771 394
R1909 VSS.n1296 VSS.n771 394
R1910 VSS.n1296 VSS.n765 394
R1911 VSS.n1304 VSS.n765 394
R1912 VSS.n1304 VSS.n763 394
R1913 VSS.n1308 VSS.n763 394
R1914 VSS.n1308 VSS.n757 394
R1915 VSS.n1316 VSS.n757 394
R1916 VSS.n1316 VSS.n755 394
R1917 VSS.n1320 VSS.n755 394
R1918 VSS.n1320 VSS.n749 394
R1919 VSS.n1329 VSS.n749 394
R1920 VSS.n1329 VSS.n747 394
R1921 VSS.n1333 VSS.n747 394
R1922 VSS.n1333 VSS.n742 394
R1923 VSS.n1342 VSS.n742 394
R1924 VSS.n1342 VSS.n740 394
R1925 VSS.n1346 VSS.n740 394
R1926 VSS.n1346 VSS.n735 394
R1927 VSS.n1355 VSS.n735 394
R1928 VSS.n1355 VSS.n733 394
R1929 VSS.n1359 VSS.n733 394
R1930 VSS.n1359 VSS.n728 394
R1931 VSS.n1369 VSS.n728 394
R1932 VSS.n1369 VSS.n726 394
R1933 VSS.n1373 VSS.n726 394
R1934 VSS.n1373 VSS.n722 394
R1935 VSS.n1788 VSS.n1616 281.082
R1936 VSS.n1978 VSS.n1977 233.52
R1937 VSS.n2335 VSS.n2334 218.815
R1938 VSS.n2335 VSS.n168 218.815
R1939 VSS.n2335 VSS.n169 218.815
R1940 VSS.n2335 VSS.n170 218.815
R1941 VSS.n2335 VSS.n171 218.815
R1942 VSS.n2335 VSS.n172 218.815
R1943 VSS.n2335 VSS.n173 218.815
R1944 VSS.n2335 VSS.n174 218.815
R1945 VSS.n2335 VSS.n175 218.815
R1946 VSS.n2335 VSS.n176 218.815
R1947 VSS.n2335 VSS.n177 218.815
R1948 VSS.n2335 VSS.n178 218.815
R1949 VSS.n2335 VSS.n179 218.815
R1950 VSS.n2335 VSS.n180 218.815
R1951 VSS.n2335 VSS.n181 218.815
R1952 VSS.n2335 VSS.n182 218.815
R1953 VSS.n2335 VSS.n183 218.815
R1954 VSS.n2335 VSS.n184 218.815
R1955 VSS.n2335 VSS.n185 218.815
R1956 VSS.n2335 VSS.n186 218.815
R1957 VSS.n1717 VSS.n1716 218.815
R1958 VSS.n1717 VSS.n1637 218.815
R1959 VSS.n1717 VSS.n1636 218.815
R1960 VSS.n1717 VSS.n1635 218.815
R1961 VSS.n1717 VSS.n1634 218.815
R1962 VSS.n1717 VSS.n1633 218.815
R1963 VSS.n1717 VSS.n1632 218.815
R1964 VSS.n1717 VSS.n1631 218.815
R1965 VSS.n1717 VSS.n1630 218.815
R1966 VSS.n1717 VSS.n1629 218.815
R1967 VSS.n1717 VSS.n1628 218.815
R1968 VSS.n1717 VSS.n1627 218.815
R1969 VSS.n1717 VSS.n1626 218.815
R1970 VSS.n1717 VSS.n1625 218.815
R1971 VSS.n1717 VSS.n1624 218.815
R1972 VSS.n1717 VSS.n1623 218.815
R1973 VSS.n1717 VSS.n1622 218.815
R1974 VSS.n1717 VSS.n1621 218.815
R1975 VSS.n1717 VSS.n1620 218.815
R1976 VSS.n1717 VSS.n1619 218.815
R1977 VSS.n1888 VSS.n1887 218.815
R1978 VSS.n1888 VSS.n1530 218.815
R1979 VSS.n2092 VSS.n2091 218.815
R1980 VSS.n2092 VSS.n678 218.815
R1981 VSS.n2092 VSS.n679 218.815
R1982 VSS.n2092 VSS.n680 218.815
R1983 VSS.n2092 VSS.n681 218.815
R1984 VSS.n2092 VSS.n682 218.815
R1985 VSS.n2092 VSS.n683 218.815
R1986 VSS.n2092 VSS.n684 218.815
R1987 VSS.n2092 VSS.n685 218.815
R1988 VSS.n2092 VSS.n686 218.815
R1989 VSS.n2092 VSS.n687 218.815
R1990 VSS.n2092 VSS.n688 218.815
R1991 VSS.n2092 VSS.n689 218.815
R1992 VSS.n2093 VSS.n2092 218.815
R1993 VSS.n1977 VSS.n1976 218.815
R1994 VSS.n1977 VSS.n1902 218.815
R1995 VSS.n1977 VSS.n1901 218.815
R1996 VSS.n1977 VSS.n1900 218.815
R1997 VSS.n1977 VSS.n1899 218.815
R1998 VSS.n1977 VSS.n1898 218.815
R1999 VSS.n1977 VSS.n1897 218.815
R2000 VSS.n1977 VSS.n1896 218.815
R2001 VSS.n1977 VSS.n1895 218.815
R2002 VSS.n1977 VSS.n1894 218.815
R2003 VSS.n1977 VSS.n1893 218.815
R2004 VSS.n1977 VSS.n1892 218.815
R2005 VSS.n1977 VSS.n1891 218.815
R2006 VSS.n1977 VSS.n1890 218.815
R2007 VSS.n1977 VSS.n1889 218.815
R2008 VSS.n2124 VSS.n2123 218.815
R2009 VSS.n2123 VSS.n321 218.815
R2010 VSS.n2123 VSS.n322 218.815
R2011 VSS.n2123 VSS.n323 218.815
R2012 VSS.n2123 VSS.n324 218.815
R2013 VSS.n2123 VSS.n325 218.815
R2014 VSS.n2123 VSS.n326 218.815
R2015 VSS.n2123 VSS.n327 218.815
R2016 VSS.n2123 VSS.n328 218.815
R2017 VSS.n2123 VSS.n329 218.815
R2018 VSS.n2123 VSS.n330 218.815
R2019 VSS.n2123 VSS.n331 218.815
R2020 VSS.n2123 VSS.n332 218.815
R2021 VSS.n2123 VSS.n333 218.815
R2022 VSS.n2123 VSS.n334 218.815
R2023 VSS.n2123 VSS.n335 218.815
R2024 VSS.n2123 VSS.n336 218.815
R2025 VSS.n2123 VSS.n337 218.815
R2026 VSS.n2123 VSS.n338 218.815
R2027 VSS.n2123 VSS.n339 218.815
R2028 VSS.n2123 VSS.n340 218.815
R2029 VSS.n2123 VSS.n341 218.815
R2030 VSS.n2123 VSS.n342 218.815
R2031 VSS.n2226 VSS.n210 218.815
R2032 VSS.n2226 VSS.n209 218.815
R2033 VSS.n2226 VSS.n208 218.815
R2034 VSS.n2226 VSS.n207 218.815
R2035 VSS.n2226 VSS.n206 218.815
R2036 VSS.n2226 VSS.n205 218.815
R2037 VSS.n2226 VSS.n204 218.815
R2038 VSS.n2226 VSS.n203 218.815
R2039 VSS.n2226 VSS.n202 218.815
R2040 VSS.n2226 VSS.n201 218.815
R2041 VSS.n2226 VSS.n200 218.815
R2042 VSS.n2226 VSS.n199 218.815
R2043 VSS.n2226 VSS.n198 218.815
R2044 VSS.n2226 VSS.n197 218.815
R2045 VSS.n2226 VSS.n196 218.815
R2046 VSS.n2226 VSS.n195 218.815
R2047 VSS.n2226 VSS.n194 218.815
R2048 VSS.n2226 VSS.n193 218.815
R2049 VSS.n2226 VSS.n192 218.815
R2050 VSS.n2226 VSS.n191 218.815
R2051 VSS.n2226 VSS.n190 218.815
R2052 VSS.n2226 VSS.n189 218.815
R2053 VSS.n2226 VSS.n188 218.815
R2054 VSS.n2107 VSS.n2106 218.815
R2055 VSS.n2107 VSS.n670 218.815
R2056 VSS.n1964 VSS.n239 218.815
R2057 VSS.n1969 VSS.n239 218.815
R2058 VSS.n1963 VSS.n239 218.815
R2059 VSS.n1496 VSS.n1495 218.815
R2060 VSS.n1496 VSS.n691 218.815
R2061 VSS.n1496 VSS.n692 218.815
R2062 VSS.n1496 VSS.n693 218.815
R2063 VSS.n1496 VSS.n694 218.815
R2064 VSS.n1496 VSS.n695 218.815
R2065 VSS.n1496 VSS.n696 218.815
R2066 VSS.n1496 VSS.n697 218.815
R2067 VSS.n1496 VSS.n698 218.815
R2068 VSS.n1496 VSS.n699 218.815
R2069 VSS.n1496 VSS.n700 218.815
R2070 VSS.n1496 VSS.n701 218.815
R2071 VSS.n1496 VSS.n702 218.815
R2072 VSS.n1496 VSS.n703 218.815
R2073 VSS.n1496 VSS.n704 218.815
R2074 VSS.n1496 VSS.n705 218.815
R2075 VSS.n1496 VSS.n706 218.815
R2076 VSS.n1496 VSS.n707 218.815
R2077 VSS.n1496 VSS.n708 218.815
R2078 VSS.n1496 VSS.n709 218.815
R2079 VSS.n1496 VSS.n710 218.815
R2080 VSS.n1496 VSS.n711 218.815
R2081 VSS.n1496 VSS.n712 218.815
R2082 VSS.n1496 VSS.n713 218.815
R2083 VSS.n1496 VSS.n714 218.815
R2084 VSS.n1496 VSS.n715 218.815
R2085 VSS.n1496 VSS.n716 218.815
R2086 VSS.n1496 VSS.n717 218.815
R2087 VSS.n1496 VSS.n718 218.815
R2088 VSS.n1103 VSS.n671 218.815
R2089 VSS.n1102 VSS.n671 218.815
R2090 VSS.n1110 VSS.n671 218.815
R2091 VSS.n867 VSS.n671 218.815
R2092 VSS.n1117 VSS.n671 218.815
R2093 VSS.n864 VSS.n671 218.815
R2094 VSS.n1124 VSS.n671 218.815
R2095 VSS.n861 VSS.n671 218.815
R2096 VSS.n1131 VSS.n671 218.815
R2097 VSS.n858 VSS.n671 218.815
R2098 VSS.n1138 VSS.n671 218.815
R2099 VSS.n855 VSS.n671 218.815
R2100 VSS.n1145 VSS.n671 218.815
R2101 VSS.n852 VSS.n671 218.815
R2102 VSS.n1152 VSS.n671 218.815
R2103 VSS.n849 VSS.n671 218.815
R2104 VSS.n1159 VSS.n671 218.815
R2105 VSS.n846 VSS.n671 218.815
R2106 VSS.n1166 VSS.n671 218.815
R2107 VSS.n843 VSS.n671 218.815
R2108 VSS.n1173 VSS.n671 218.815
R2109 VSS.n840 VSS.n671 218.815
R2110 VSS.n1180 VSS.n671 218.815
R2111 VSS.n837 VSS.n671 218.815
R2112 VSS.n1187 VSS.n671 218.815
R2113 VSS.n834 VSS.n671 218.815
R2114 VSS.n1194 VSS.n671 218.815
R2115 VSS.n831 VSS.n671 218.815
R2116 VSS.n1201 VSS.n671 218.815
R2117 VSS.n828 VSS.n671 218.815
R2118 VSS.n2092 VSS.n677 210.695
R2119 VSS.n503 VSS.n188 147.374
R2120 VSS.n507 VSS.n189 147.374
R2121 VSS.n511 VSS.n190 147.374
R2122 VSS.n515 VSS.n191 147.374
R2123 VSS.n519 VSS.n192 147.374
R2124 VSS.n523 VSS.n193 147.374
R2125 VSS.n527 VSS.n194 147.374
R2126 VSS.n531 VSS.n195 147.374
R2127 VSS.n535 VSS.n196 147.374
R2128 VSS.n539 VSS.n197 147.374
R2129 VSS.n543 VSS.n198 147.374
R2130 VSS.n547 VSS.n199 147.374
R2131 VSS.n551 VSS.n200 147.374
R2132 VSS.n555 VSS.n201 147.374
R2133 VSS.n559 VSS.n202 147.374
R2134 VSS.n563 VSS.n203 147.374
R2135 VSS.n567 VSS.n204 147.374
R2136 VSS.n571 VSS.n205 147.374
R2137 VSS.n575 VSS.n206 147.374
R2138 VSS.n579 VSS.n207 147.374
R2139 VSS.n583 VSS.n208 147.374
R2140 VSS.n587 VSS.n209 147.374
R2141 VSS.n590 VSS.n210 147.374
R2142 VSS.n2124 VSS.n317 147.374
R2143 VSS.n344 VSS.n321 147.374
R2144 VSS.n348 VSS.n322 147.374
R2145 VSS.n352 VSS.n323 147.374
R2146 VSS.n356 VSS.n324 147.374
R2147 VSS.n360 VSS.n325 147.374
R2148 VSS.n364 VSS.n326 147.374
R2149 VSS.n368 VSS.n327 147.374
R2150 VSS.n372 VSS.n328 147.374
R2151 VSS.n376 VSS.n329 147.374
R2152 VSS.n380 VSS.n330 147.374
R2153 VSS.n384 VSS.n331 147.374
R2154 VSS.n388 VSS.n332 147.374
R2155 VSS.n392 VSS.n333 147.374
R2156 VSS.n396 VSS.n334 147.374
R2157 VSS.n400 VSS.n335 147.374
R2158 VSS.n404 VSS.n336 147.374
R2159 VSS.n408 VSS.n337 147.374
R2160 VSS.n412 VSS.n338 147.374
R2161 VSS.n416 VSS.n339 147.374
R2162 VSS.n420 VSS.n340 147.374
R2163 VSS.n424 VSS.n341 147.374
R2164 VSS.n428 VSS.n342 147.374
R2165 VSS.n1908 VSS.n1889 147.374
R2166 VSS.n1912 VSS.n1890 147.374
R2167 VSS.n1916 VSS.n1891 147.374
R2168 VSS.n1920 VSS.n1892 147.374
R2169 VSS.n1924 VSS.n1893 147.374
R2170 VSS.n1928 VSS.n1894 147.374
R2171 VSS.n1932 VSS.n1895 147.374
R2172 VSS.n1936 VSS.n1896 147.374
R2173 VSS.n1940 VSS.n1897 147.374
R2174 VSS.n1944 VSS.n1898 147.374
R2175 VSS.n1948 VSS.n1899 147.374
R2176 VSS.n1952 VSS.n1900 147.374
R2177 VSS.n1956 VSS.n1901 147.374
R2178 VSS.n1959 VSS.n1902 147.374
R2179 VSS.n1976 VSS.n1975 147.374
R2180 VSS.n1971 VSS.n1963 147.374
R2181 VSS.n1969 VSS.n1968 147.374
R2182 VSS.n1964 VSS.n243 147.374
R2183 VSS.n2091 VSS.n2090 147.374
R2184 VSS.n2085 VSS.n678 147.374
R2185 VSS.n2082 VSS.n679 147.374
R2186 VSS.n2078 VSS.n680 147.374
R2187 VSS.n2074 VSS.n681 147.374
R2188 VSS.n2070 VSS.n682 147.374
R2189 VSS.n2066 VSS.n683 147.374
R2190 VSS.n2062 VSS.n684 147.374
R2191 VSS.n2058 VSS.n685 147.374
R2192 VSS.n2054 VSS.n686 147.374
R2193 VSS.n2050 VSS.n687 147.374
R2194 VSS.n2046 VSS.n688 147.374
R2195 VSS.n2042 VSS.n689 147.374
R2196 VSS.n2093 VSS.n676 147.374
R2197 VSS.n2106 VSS.n2105 147.374
R2198 VSS.n2100 VSS.n670 147.374
R2199 VSS.n1887 VSS.n1886 147.374
R2200 VSS.n1881 VSS.n1530 147.374
R2201 VSS.n1642 VSS.n1619 147.374
R2202 VSS.n1646 VSS.n1620 147.374
R2203 VSS.n1650 VSS.n1621 147.374
R2204 VSS.n1654 VSS.n1622 147.374
R2205 VSS.n1658 VSS.n1623 147.374
R2206 VSS.n1662 VSS.n1624 147.374
R2207 VSS.n1666 VSS.n1625 147.374
R2208 VSS.n1670 VSS.n1626 147.374
R2209 VSS.n1674 VSS.n1627 147.374
R2210 VSS.n1678 VSS.n1628 147.374
R2211 VSS.n1682 VSS.n1629 147.374
R2212 VSS.n1686 VSS.n1630 147.374
R2213 VSS.n1690 VSS.n1631 147.374
R2214 VSS.n1694 VSS.n1632 147.374
R2215 VSS.n1698 VSS.n1633 147.374
R2216 VSS.n1702 VSS.n1634 147.374
R2217 VSS.n1706 VSS.n1635 147.374
R2218 VSS.n1710 VSS.n1636 147.374
R2219 VSS.n1638 VSS.n1637 147.374
R2220 VSS.n1716 VSS.n123 147.374
R2221 VSS.n2334 VSS.n165 147.374
R2222 VSS.n2329 VSS.n168 147.374
R2223 VSS.n2326 VSS.n169 147.374
R2224 VSS.n2322 VSS.n170 147.374
R2225 VSS.n2318 VSS.n171 147.374
R2226 VSS.n2314 VSS.n172 147.374
R2227 VSS.n2310 VSS.n173 147.374
R2228 VSS.n2306 VSS.n174 147.374
R2229 VSS.n2302 VSS.n175 147.374
R2230 VSS.n2298 VSS.n176 147.374
R2231 VSS.n2294 VSS.n177 147.374
R2232 VSS.n2290 VSS.n178 147.374
R2233 VSS.n2286 VSS.n179 147.374
R2234 VSS.n2282 VSS.n180 147.374
R2235 VSS.n2278 VSS.n181 147.374
R2236 VSS.n2274 VSS.n182 147.374
R2237 VSS.n2270 VSS.n183 147.374
R2238 VSS.n2266 VSS.n184 147.374
R2239 VSS.n2262 VSS.n185 147.374
R2240 VSS.n2258 VSS.n186 147.374
R2241 VSS.n2334 VSS.n2333 147.374
R2242 VSS.n2327 VSS.n168 147.374
R2243 VSS.n2323 VSS.n169 147.374
R2244 VSS.n2319 VSS.n170 147.374
R2245 VSS.n2315 VSS.n171 147.374
R2246 VSS.n2311 VSS.n172 147.374
R2247 VSS.n2307 VSS.n173 147.374
R2248 VSS.n2303 VSS.n174 147.374
R2249 VSS.n2299 VSS.n175 147.374
R2250 VSS.n2295 VSS.n176 147.374
R2251 VSS.n2291 VSS.n177 147.374
R2252 VSS.n2287 VSS.n178 147.374
R2253 VSS.n2283 VSS.n179 147.374
R2254 VSS.n2279 VSS.n180 147.374
R2255 VSS.n2275 VSS.n181 147.374
R2256 VSS.n2271 VSS.n182 147.374
R2257 VSS.n2267 VSS.n183 147.374
R2258 VSS.n2263 VSS.n184 147.374
R2259 VSS.n2259 VSS.n185 147.374
R2260 VSS.n2255 VSS.n186 147.374
R2261 VSS.n1716 VSS.n1715 147.374
R2262 VSS.n1711 VSS.n1637 147.374
R2263 VSS.n1707 VSS.n1636 147.374
R2264 VSS.n1703 VSS.n1635 147.374
R2265 VSS.n1699 VSS.n1634 147.374
R2266 VSS.n1695 VSS.n1633 147.374
R2267 VSS.n1691 VSS.n1632 147.374
R2268 VSS.n1687 VSS.n1631 147.374
R2269 VSS.n1683 VSS.n1630 147.374
R2270 VSS.n1679 VSS.n1629 147.374
R2271 VSS.n1675 VSS.n1628 147.374
R2272 VSS.n1671 VSS.n1627 147.374
R2273 VSS.n1667 VSS.n1626 147.374
R2274 VSS.n1663 VSS.n1625 147.374
R2275 VSS.n1659 VSS.n1624 147.374
R2276 VSS.n1655 VSS.n1623 147.374
R2277 VSS.n1651 VSS.n1622 147.374
R2278 VSS.n1647 VSS.n1621 147.374
R2279 VSS.n1643 VSS.n1620 147.374
R2280 VSS.n1639 VSS.n1619 147.374
R2281 VSS.n1887 VSS.n1533 147.374
R2282 VSS.n1879 VSS.n1530 147.374
R2283 VSS.n2091 VSS.n1498 147.374
R2284 VSS.n2083 VSS.n678 147.374
R2285 VSS.n2079 VSS.n679 147.374
R2286 VSS.n2075 VSS.n680 147.374
R2287 VSS.n2071 VSS.n681 147.374
R2288 VSS.n2067 VSS.n682 147.374
R2289 VSS.n2063 VSS.n683 147.374
R2290 VSS.n2059 VSS.n684 147.374
R2291 VSS.n2055 VSS.n685 147.374
R2292 VSS.n2051 VSS.n686 147.374
R2293 VSS.n2047 VSS.n687 147.374
R2294 VSS.n2043 VSS.n688 147.374
R2295 VSS.n2039 VSS.n689 147.374
R2296 VSS.n2094 VSS.n2093 147.374
R2297 VSS.n1976 VSS.n1903 147.374
R2298 VSS.n1957 VSS.n1902 147.374
R2299 VSS.n1953 VSS.n1901 147.374
R2300 VSS.n1949 VSS.n1900 147.374
R2301 VSS.n1945 VSS.n1899 147.374
R2302 VSS.n1941 VSS.n1898 147.374
R2303 VSS.n1937 VSS.n1897 147.374
R2304 VSS.n1933 VSS.n1896 147.374
R2305 VSS.n1929 VSS.n1895 147.374
R2306 VSS.n1925 VSS.n1894 147.374
R2307 VSS.n1921 VSS.n1893 147.374
R2308 VSS.n1917 VSS.n1892 147.374
R2309 VSS.n1913 VSS.n1891 147.374
R2310 VSS.n1909 VSS.n1890 147.374
R2311 VSS.n1905 VSS.n1889 147.374
R2312 VSS.n2125 VSS.n2124 147.374
R2313 VSS.n347 VSS.n321 147.374
R2314 VSS.n351 VSS.n322 147.374
R2315 VSS.n355 VSS.n323 147.374
R2316 VSS.n359 VSS.n324 147.374
R2317 VSS.n363 VSS.n325 147.374
R2318 VSS.n367 VSS.n326 147.374
R2319 VSS.n371 VSS.n327 147.374
R2320 VSS.n375 VSS.n328 147.374
R2321 VSS.n379 VSS.n329 147.374
R2322 VSS.n383 VSS.n330 147.374
R2323 VSS.n387 VSS.n331 147.374
R2324 VSS.n391 VSS.n332 147.374
R2325 VSS.n395 VSS.n333 147.374
R2326 VSS.n399 VSS.n334 147.374
R2327 VSS.n403 VSS.n335 147.374
R2328 VSS.n407 VSS.n336 147.374
R2329 VSS.n411 VSS.n337 147.374
R2330 VSS.n415 VSS.n338 147.374
R2331 VSS.n419 VSS.n339 147.374
R2332 VSS.n423 VSS.n340 147.374
R2333 VSS.n427 VSS.n341 147.374
R2334 VSS.n343 VSS.n342 147.374
R2335 VSS.n588 VSS.n210 147.374
R2336 VSS.n584 VSS.n209 147.374
R2337 VSS.n580 VSS.n208 147.374
R2338 VSS.n576 VSS.n207 147.374
R2339 VSS.n572 VSS.n206 147.374
R2340 VSS.n568 VSS.n205 147.374
R2341 VSS.n564 VSS.n204 147.374
R2342 VSS.n560 VSS.n203 147.374
R2343 VSS.n556 VSS.n202 147.374
R2344 VSS.n552 VSS.n201 147.374
R2345 VSS.n548 VSS.n200 147.374
R2346 VSS.n544 VSS.n199 147.374
R2347 VSS.n540 VSS.n198 147.374
R2348 VSS.n536 VSS.n197 147.374
R2349 VSS.n532 VSS.n196 147.374
R2350 VSS.n528 VSS.n195 147.374
R2351 VSS.n524 VSS.n194 147.374
R2352 VSS.n520 VSS.n193 147.374
R2353 VSS.n516 VSS.n192 147.374
R2354 VSS.n512 VSS.n191 147.374
R2355 VSS.n508 VSS.n190 147.374
R2356 VSS.n504 VSS.n189 147.374
R2357 VSS.n213 VSS.n188 147.374
R2358 VSS.n2106 VSS.n673 147.374
R2359 VSS.n2098 VSS.n670 147.374
R2360 VSS.n1965 VSS.n1964 147.374
R2361 VSS.n1970 VSS.n1969 147.374
R2362 VSS.n1963 VSS.n1904 147.374
R2363 VSS.n1495 VSS.n1494 147.374
R2364 VSS.n1489 VSS.n691 147.374
R2365 VSS.n1486 VSS.n692 147.374
R2366 VSS.n1482 VSS.n693 147.374
R2367 VSS.n1478 VSS.n694 147.374
R2368 VSS.n1474 VSS.n695 147.374
R2369 VSS.n1470 VSS.n696 147.374
R2370 VSS.n1466 VSS.n697 147.374
R2371 VSS.n1462 VSS.n698 147.374
R2372 VSS.n1458 VSS.n699 147.374
R2373 VSS.n1454 VSS.n700 147.374
R2374 VSS.n1450 VSS.n701 147.374
R2375 VSS.n1446 VSS.n702 147.374
R2376 VSS.n1442 VSS.n703 147.374
R2377 VSS.n1438 VSS.n704 147.374
R2378 VSS.n1434 VSS.n705 147.374
R2379 VSS.n1430 VSS.n706 147.374
R2380 VSS.n1426 VSS.n707 147.374
R2381 VSS.n1422 VSS.n708 147.374
R2382 VSS.n1418 VSS.n709 147.374
R2383 VSS.n1414 VSS.n710 147.374
R2384 VSS.n1410 VSS.n711 147.374
R2385 VSS.n1406 VSS.n712 147.374
R2386 VSS.n1402 VSS.n713 147.374
R2387 VSS.n1398 VSS.n714 147.374
R2388 VSS.n1394 VSS.n715 147.374
R2389 VSS.n1390 VSS.n716 147.374
R2390 VSS.n1386 VSS.n717 147.374
R2391 VSS.n1382 VSS.n718 147.374
R2392 VSS.n1203 VSS.n828 147.374
R2393 VSS.n1201 VSS.n1200 147.374
R2394 VSS.n1196 VSS.n831 147.374
R2395 VSS.n1194 VSS.n1193 147.374
R2396 VSS.n1189 VSS.n834 147.374
R2397 VSS.n1187 VSS.n1186 147.374
R2398 VSS.n1182 VSS.n837 147.374
R2399 VSS.n1180 VSS.n1179 147.374
R2400 VSS.n1175 VSS.n840 147.374
R2401 VSS.n1173 VSS.n1172 147.374
R2402 VSS.n1168 VSS.n843 147.374
R2403 VSS.n1166 VSS.n1165 147.374
R2404 VSS.n1161 VSS.n846 147.374
R2405 VSS.n1159 VSS.n1158 147.374
R2406 VSS.n1154 VSS.n849 147.374
R2407 VSS.n1152 VSS.n1151 147.374
R2408 VSS.n1147 VSS.n852 147.374
R2409 VSS.n1145 VSS.n1144 147.374
R2410 VSS.n1140 VSS.n855 147.374
R2411 VSS.n1138 VSS.n1137 147.374
R2412 VSS.n1133 VSS.n858 147.374
R2413 VSS.n1131 VSS.n1130 147.374
R2414 VSS.n1126 VSS.n861 147.374
R2415 VSS.n1124 VSS.n1123 147.374
R2416 VSS.n1119 VSS.n864 147.374
R2417 VSS.n1117 VSS.n1116 147.374
R2418 VSS.n1112 VSS.n867 147.374
R2419 VSS.n1110 VSS.n1109 147.374
R2420 VSS.n1105 VSS.n1102 147.374
R2421 VSS.n1103 VSS.n825 147.374
R2422 VSS.n1495 VSS.n721 147.374
R2423 VSS.n1487 VSS.n691 147.374
R2424 VSS.n1483 VSS.n692 147.374
R2425 VSS.n1479 VSS.n693 147.374
R2426 VSS.n1475 VSS.n694 147.374
R2427 VSS.n1471 VSS.n695 147.374
R2428 VSS.n1467 VSS.n696 147.374
R2429 VSS.n1463 VSS.n697 147.374
R2430 VSS.n1459 VSS.n698 147.374
R2431 VSS.n1455 VSS.n699 147.374
R2432 VSS.n1451 VSS.n700 147.374
R2433 VSS.n1447 VSS.n701 147.374
R2434 VSS.n1443 VSS.n702 147.374
R2435 VSS.n1439 VSS.n703 147.374
R2436 VSS.n1435 VSS.n704 147.374
R2437 VSS.n1431 VSS.n705 147.374
R2438 VSS.n1427 VSS.n706 147.374
R2439 VSS.n1423 VSS.n707 147.374
R2440 VSS.n1419 VSS.n708 147.374
R2441 VSS.n1415 VSS.n709 147.374
R2442 VSS.n1411 VSS.n710 147.374
R2443 VSS.n1407 VSS.n711 147.374
R2444 VSS.n1403 VSS.n712 147.374
R2445 VSS.n1399 VSS.n713 147.374
R2446 VSS.n1395 VSS.n714 147.374
R2447 VSS.n1391 VSS.n715 147.374
R2448 VSS.n1387 VSS.n716 147.374
R2449 VSS.n1383 VSS.n717 147.374
R2450 VSS.n1379 VSS.n718 147.374
R2451 VSS.n1104 VSS.n1103 147.374
R2452 VSS.n1102 VSS.n868 147.374
R2453 VSS.n1111 VSS.n1110 147.374
R2454 VSS.n867 VSS.n865 147.374
R2455 VSS.n1118 VSS.n1117 147.374
R2456 VSS.n864 VSS.n862 147.374
R2457 VSS.n1125 VSS.n1124 147.374
R2458 VSS.n861 VSS.n859 147.374
R2459 VSS.n1132 VSS.n1131 147.374
R2460 VSS.n858 VSS.n856 147.374
R2461 VSS.n1139 VSS.n1138 147.374
R2462 VSS.n855 VSS.n853 147.374
R2463 VSS.n1146 VSS.n1145 147.374
R2464 VSS.n852 VSS.n850 147.374
R2465 VSS.n1153 VSS.n1152 147.374
R2466 VSS.n849 VSS.n847 147.374
R2467 VSS.n1160 VSS.n1159 147.374
R2468 VSS.n846 VSS.n844 147.374
R2469 VSS.n1167 VSS.n1166 147.374
R2470 VSS.n843 VSS.n841 147.374
R2471 VSS.n1174 VSS.n1173 147.374
R2472 VSS.n840 VSS.n838 147.374
R2473 VSS.n1181 VSS.n1180 147.374
R2474 VSS.n837 VSS.n835 147.374
R2475 VSS.n1188 VSS.n1187 147.374
R2476 VSS.n834 VSS.n832 147.374
R2477 VSS.n1195 VSS.n1194 147.374
R2478 VSS.n831 VSS.n829 147.374
R2479 VSS.n1202 VSS.n1201 147.374
R2480 VSS.n828 VSS.n826 147.374
R2481 VSS.n1979 VSS.n1978 119.394
R2482 VSS.n1985 VSS.n1526 119.394
R2483 VSS.n1986 VSS.n1985 119.394
R2484 VSS.n1987 VSS.n1986 119.394
R2485 VSS.n1993 VSS.n1522 119.394
R2486 VSS.n1994 VSS.n1993 119.394
R2487 VSS.n1995 VSS.n1994 119.394
R2488 VSS.n2001 VSS.n1518 119.394
R2489 VSS.n2002 VSS.n2001 119.394
R2490 VSS.n2003 VSS.n2002 119.394
R2491 VSS.n2009 VSS.n1514 119.394
R2492 VSS.n2010 VSS.n2009 119.394
R2493 VSS.n2011 VSS.n1510 119.394
R2494 VSS.n2017 VSS.n1510 119.394
R2495 VSS.n2018 VSS.n2017 119.394
R2496 VSS.n2025 VSS.n1506 119.394
R2497 VSS.n2026 VSS.n2025 119.394
R2498 VSS.n2027 VSS.n1502 119.394
R2499 VSS.n2033 VSS.n1502 119.394
R2500 VSS.n2034 VSS.n2033 119.394
R2501 VSS.n2035 VSS.n677 119.394
R2502 VSS.t4 VSS.n1514 117.638
R2503 VSS.t53 VSS.n484 114.742
R2504 VSS.n485 VSS.t53 114.742
R2505 VSS.t145 VSS.n486 114.742
R2506 VSS.n487 VSS.t145 114.742
R2507 VSS.t50 VSS.n488 114.742
R2508 VSS.n489 VSS.t50 114.742
R2509 VSS.t140 VSS.n490 114.742
R2510 VSS.n491 VSS.t140 114.742
R2511 VSS.t170 VSS.n492 114.742
R2512 VSS.n493 VSS.t170 114.742
R2513 VSS.t91 VSS.n494 114.742
R2514 VSS.n495 VSS.t91 114.742
R2515 VSS.t131 VSS.n496 114.742
R2516 VSS.n497 VSS.t131 114.742
R2517 VSS.t199 VSS.n462 114.742
R2518 VSS.t107 VSS.n464 114.742
R2519 VSS.t195 VSS.n466 114.742
R2520 VSS.t105 VSS.n468 114.742
R2521 VSS.t127 VSS.n470 114.742
R2522 VSS.t26 VSS.n472 114.742
R2523 VSS.t93 VSS.n474 114.742
R2524 VSS.n907 VSS.t47 114.742
R2525 VSS.n914 VSS.t83 114.742
R2526 VSS.t179 VSS.n927 114.742
R2527 VSS.t205 VSS.n929 114.742
R2528 VSS.t123 VSS.n931 114.742
R2529 VSS.t63 VSS.n933 114.742
R2530 VSS.t207 VSS.n935 114.742
R2531 VSS.n940 VSS.t71 114.742
R2532 VSS.t109 VSS.n941 114.742
R2533 VSS.n942 VSS.t109 114.742
R2534 VSS.t60 VSS.n943 114.742
R2535 VSS.n944 VSS.t60 114.742
R2536 VSS.t153 VSS.n945 114.742
R2537 VSS.n946 VSS.t153 114.742
R2538 VSS.t125 VSS.n947 114.742
R2539 VSS.n948 VSS.t125 114.742
R2540 VSS.t101 VSS.n949 114.742
R2541 VSS.n102 VSS.t97 114.742
R2542 VSS.n66 VSS.t33 114.742
R2543 VSS.t33 VSS.n65 114.742
R2544 VSS.n1077 VSS.t136 114.742
R2545 VSS.t136 VSS.n1076 114.742
R2546 VSS.n1075 VSS.t37 114.742
R2547 VSS.t37 VSS.n1074 114.742
R2548 VSS.n1073 VSS.t138 114.742
R2549 VSS.t138 VSS.n1072 114.742
R2550 VSS.n1071 VSS.t40 114.742
R2551 VSS.t40 VSS.n1070 114.742
R2552 VSS.n1069 VSS.t193 114.742
R2553 VSS.t193 VSS.n1068 114.742
R2554 VSS.n1067 VSS.t113 114.742
R2555 VSS.t113 VSS.n1066 114.742
R2556 VSS.n1065 VSS.t66 114.742
R2557 VSS.t66 VSS.n1064 114.742
R2558 VSS.n1041 VSS.t164 114.742
R2559 VSS.n1039 VSS.t79 114.742
R2560 VSS.n1037 VSS.t121 114.742
R2561 VSS.n1035 VSS.t201 114.742
R2562 VSS.n1033 VSS.t58 114.742
R2563 VSS.n1031 VSS.t151 114.742
R2564 VSS.n1029 VSS.t55 114.742
R2565 VSS.n463 VSS.t199 114.742
R2566 VSS.n465 VSS.t107 114.742
R2567 VSS.n467 VSS.t195 114.742
R2568 VSS.n469 VSS.t105 114.742
R2569 VSS.n471 VSS.t127 114.742
R2570 VSS.n473 VSS.t26 114.742
R2571 VSS.n475 VSS.t93 114.742
R2572 VSS.n917 VSS.t88 114.742
R2573 VSS.n924 VSS.t155 114.742
R2574 VSS.n926 VSS.t161 114.742
R2575 VSS.n928 VSS.t179 114.742
R2576 VSS.n930 VSS.t205 114.742
R2577 VSS.n932 VSS.t123 114.742
R2578 VSS.n934 VSS.t63 114.742
R2579 VSS.t97 VSS.n101 114.742
R2580 VSS.t81 VSS.n1042 114.742
R2581 VSS.t164 VSS.n1040 114.742
R2582 VSS.t79 VSS.n1038 114.742
R2583 VSS.t121 VSS.n1036 114.742
R2584 VSS.t201 VSS.n1034 114.742
R2585 VSS.t58 VSS.n1032 114.742
R2586 VSS.t151 VSS.n1030 114.742
R2587 VSS.t55 VSS.n1028 114.742
R2588 VSS.n1022 VSS.t35 114.707
R2589 VSS.n1021 VSS.t175 114.707
R2590 VSS.n1048 VSS.t203 114.707
R2591 VSS.n995 VSS.t74 114.707
R2592 VSS.n973 VSS.t111 114.707
R2593 VSS.n971 VSS.t24 114.707
R2594 VSS.n971 VSS.t95 114.707
R2595 VSS.n1002 VSS.t115 114.707
R2596 VSS.n967 VSS.t44 114.397
R2597 VSS.n1020 VSS.t181 114.397
R2598 VSS.n1052 VSS.t129 114.397
R2599 VSS.n1051 VSS.t168 114.397
R2600 VSS.n1049 VSS.t166 114.397
R2601 VSS.n994 VSS.t76 114.397
R2602 VSS.n974 VSS.t117 114.397
R2603 VSS.n1003 VSS.t119 114.397
R2604 VSS.t161 VSS.n925 114.391
R2605 VSS.n936 VSS.t207 114.391
R2606 VSS.t71 VSS.n939 114.391
R2607 VSS.n950 VSS.t101 114.391
R2608 VSS.t209 VSS.n52 114.391
R2609 VSS.n53 VSS.t209 114.391
R2610 VSS.t172 VSS.n57 114.391
R2611 VSS.n58 VSS.t172 114.391
R2612 VSS.t142 VSS.n68 114.391
R2613 VSS.n69 VSS.t142 114.391
R2614 VSS.t29 VSS.n72 114.391
R2615 VSS.n73 VSS.t29 114.391
R2616 VSS.n24 VSS.t99 114.391
R2617 VSS.t99 VSS.n22 114.391
R2618 VSS.t191 VSS.n98 114.391
R2619 VSS.n99 VSS.t191 114.391
R2620 VSS.t177 VSS.n106 114.391
R2621 VSS.n107 VSS.t177 114.391
R2622 VSS.n14 VSS.t21 114.391
R2623 VSS.t21 VSS.n12 114.391
R2624 VSS.t86 VSS.n118 114.391
R2625 VSS.n119 VSS.t86 114.391
R2626 VSS.n89 VSS.t42 114.391
R2627 VSS.t42 VSS.n88 114.391
R2628 VSS.n76 VSS.t183 114.391
R2629 VSS.t183 VSS.n29 114.391
R2630 VSS.n61 VSS.t133 114.391
R2631 VSS.t133 VSS.n41 114.391
R2632 VSS.n1096 VSS.t197 114.391
R2633 VSS.t197 VSS.n1095 114.391
R2634 VSS.t158 VSS.n1061 114.391
R2635 VSS.n1062 VSS.t158 114.391
R2636 VSS.t188 VSS.n1079 114.391
R2637 VSS.n1080 VSS.t188 114.391
R2638 VSS.n1058 VSS.t68 114.391
R2639 VSS.t68 VSS.n1057 114.391
R2640 VSS.n1043 VSS.t81 114.391
R2641 VSS.n1016 VSS.t149 114.391
R2642 VSS.t149 VSS.n1015 114.391
R2643 VSS.n1888 VSS.n1531 112.442
R2644 VSS.t2 VSS.n2010 96.5687
R2645 VSS.n2035 VSS.t61 96.5687
R2646 VSS.t3 VSS.n1518 93.0572
R2647 VSS.n1378 VSS.n1377 92.2358
R2648 VSS.n1212 VSS.n824 90.7299
R2649 VSS.n2191 VSS.n245 89.977
R2650 VSS.n483 VSS.t187 87.2694
R2651 VSS.n461 VSS.t148 87.2694
R2652 VSS.t198 VSS.n962 87.0902
R2653 VSS.n476 VSS.t132 87.0895
R2654 VSS.n477 VSS.t92 87.0895
R2655 VSS.n478 VSS.t171 87.0895
R2656 VSS.n479 VSS.t141 87.0895
R2657 VSS.n480 VSS.t52 87.0895
R2658 VSS.n481 VSS.t146 87.0895
R2659 VSS.n482 VSS.t54 87.0895
R2660 VSS.n454 VSS.t94 87.0895
R2661 VSS.n455 VSS.t28 87.0895
R2662 VSS.n456 VSS.t128 87.0895
R2663 VSS.n457 VSS.t106 87.0895
R2664 VSS.n458 VSS.t196 87.0895
R2665 VSS.n459 VSS.t108 87.0895
R2666 VSS.n460 VSS.t200 87.0895
R2667 VSS.n905 VSS.t104 87.0895
R2668 VSS.n908 VSS.t126 87.0895
R2669 VSS.n909 VSS.t154 87.0895
R2670 VSS.n910 VSS.t62 87.0895
R2671 VSS.n911 VSS.t110 87.0895
R2672 VSS.n912 VSS.t73 87.0895
R2673 VSS.t163 VSS.n922 87.0895
R2674 VSS.n921 VSS.t180 87.0895
R2675 VSS.n920 VSS.t206 87.0895
R2676 VSS.n919 VSS.t124 87.0895
R2677 VSS.n918 VSS.t65 87.0895
R2678 VSS.t208 VSS.n915 87.0895
R2679 VSS.n54 VSS.t211 87.0895
R2680 VSS.n48 VSS.t174 87.0895
R2681 VSS.n63 VSS.t135 87.0895
R2682 VSS.n40 VSS.t34 87.0895
R2683 VSS.n36 VSS.t144 87.0895
R2684 VSS.n32 VSS.t32 87.0895
R2685 VSS.t87 VSS.n10 87.0895
R2686 VSS.t23 VSS.n111 87.0895
R2687 VSS.t178 VSS.n15 87.0895
R2688 VSS.n17 VSS.t98 87.0895
R2689 VSS.t192 VSS.n18 87.0895
R2690 VSS.t100 VSS.n93 87.0895
R2691 VSS.t43 VSS.n25 87.0895
R2692 VSS.n31 VSS.t185 87.0895
R2693 VSS.n1026 VSS.t150 87.0895
R2694 VSS.n1014 VSS.t57 87.0895
R2695 VSS.n1013 VSS.t152 87.0895
R2696 VSS.n1012 VSS.t59 87.0895
R2697 VSS.n1011 VSS.t202 87.0895
R2698 VSS.n1010 VSS.t122 87.0895
R2699 VSS.n1009 VSS.t80 87.0895
R2700 VSS.n1008 VSS.t165 87.0895
R2701 VSS.n1007 VSS.t82 87.0895
R2702 VSS.n977 VSS.t190 87.0895
R2703 VSS.n978 VSS.t137 87.0895
R2704 VSS.n979 VSS.t39 87.0895
R2705 VSS.n980 VSS.t139 87.0895
R2706 VSS.n981 VSS.t41 87.0895
R2707 VSS.n982 VSS.t194 87.0895
R2708 VSS.n983 VSS.t114 87.0895
R2709 VSS.n984 VSS.t67 87.0895
R2710 VSS.n985 VSS.t160 87.0895
R2711 VSS.n988 VSS.t70 87.0895
R2712 VSS.n2128 VSS.n2127 84.7064
R2713 VSS.n660 VSS.n659 84.7064
R2714 VSS.n2338 VSS.n164 84.7064
R2715 VSS.n1493 VSS.n723 84.7064
R2716 VSS.n1906 VSS.n1528 82.0711
R2717 VSS.n2254 VSS.n2253 80.9417
R2718 VSS.n2385 VSS.n121 78.6829
R2719 VSS.n2223 VSS.n215 78.6829
R2720 VSS.n592 VSS.n591 78.6829
R2721 VSS.n1206 VSS.n1205 78.6829
R2722 VSS.n1876 VSS.n1531 77.2333
R2723 VSS.n1876 VSS.n1539 77.2333
R2724 VSS.n1870 VSS.n1539 77.2333
R2725 VSS.n1870 VSS.n1869 77.2333
R2726 VSS.n1869 VSS.n1868 77.2333
R2727 VSS.n1868 VSS.n1546 77.2333
R2728 VSS.n1862 VSS.n1546 77.2333
R2729 VSS.n1862 VSS.n1861 77.2333
R2730 VSS.n1861 VSS.n1860 77.2333
R2731 VSS.n1860 VSS.n1553 77.2333
R2732 VSS.n1854 VSS.n1553 77.2333
R2733 VSS.n1854 VSS.n1853 77.2333
R2734 VSS.n1853 VSS.n1852 77.2333
R2735 VSS.n1852 VSS.n1560 77.2333
R2736 VSS.n1846 VSS.n1560 77.2333
R2737 VSS.n1846 VSS.n1845 77.2333
R2738 VSS.n1845 VSS.n1844 77.2333
R2739 VSS.n1844 VSS.n1567 77.2333
R2740 VSS.n1838 VSS.n1567 77.2333
R2741 VSS.n1838 VSS.n1837 77.2333
R2742 VSS.n1837 VSS.n1836 77.2333
R2743 VSS.n1836 VSS.n1574 77.2333
R2744 VSS.n1830 VSS.n1829 77.2333
R2745 VSS.n1829 VSS.n1828 77.2333
R2746 VSS.n1828 VSS.n1581 77.2333
R2747 VSS.n1822 VSS.n1581 77.2333
R2748 VSS.n1822 VSS.n1821 77.2333
R2749 VSS.n1821 VSS.n1820 77.2333
R2750 VSS.n1820 VSS.n1588 77.2333
R2751 VSS.n1814 VSS.n1588 77.2333
R2752 VSS.n1814 VSS.n1813 77.2333
R2753 VSS.n1813 VSS.n1812 77.2333
R2754 VSS.n1812 VSS.n1595 77.2333
R2755 VSS.n1806 VSS.n1595 77.2333
R2756 VSS.n1806 VSS.n1805 77.2333
R2757 VSS.n1805 VSS.n1804 77.2333
R2758 VSS.n1804 VSS.n1602 77.2333
R2759 VSS.n1798 VSS.n1602 77.2333
R2760 VSS.n1798 VSS.n1797 77.2333
R2761 VSS.n1797 VSS.n1796 77.2333
R2762 VSS.n1796 VSS.n1609 77.2333
R2763 VSS.n1790 VSS.n1609 77.2333
R2764 VSS.n1790 VSS.n1789 77.2333
R2765 VSS.n1789 VSS.n1788 77.2333
R2766 VSS.n2089 VSS.n2038 77.177
R2767 VSS.n433 VSS.n431 76.1488
R2768 VSS.n436 VSS.n434 76.1488
R2769 VSS.n440 VSS.n438 76.1488
R2770 VSS.n444 VSS.n442 76.1488
R2771 VSS.n448 VSS.n446 76.1488
R2772 VSS.n452 VSS.n450 76.1488
R2773 VSS.n871 VSS.n869 76.1488
R2774 VSS.n874 VSS.n872 76.1488
R2775 VSS.n879 VSS.n877 76.1488
R2776 VSS.n884 VSS.n882 76.1488
R2777 VSS.n889 VSS.n887 76.1488
R2778 VSS.n894 VSS.n892 76.1488
R2779 VSS.n899 VSS.n897 76.1488
R2780 VSS.n904 VSS.n902 76.1488
R2781 VSS.n1979 VSS.t64 75.4993
R2782 VSS.n433 VSS.n432 75.4751
R2783 VSS.n436 VSS.n435 75.4751
R2784 VSS.n440 VSS.n439 75.4751
R2785 VSS.n444 VSS.n443 75.4751
R2786 VSS.n448 VSS.n447 75.4751
R2787 VSS.n452 VSS.n451 75.4751
R2788 VSS.n871 VSS.n870 75.4751
R2789 VSS.n874 VSS.n873 75.4751
R2790 VSS.n876 VSS.n875 75.4751
R2791 VSS.n879 VSS.n878 75.4751
R2792 VSS.n881 VSS.n880 75.4751
R2793 VSS.n884 VSS.n883 75.4751
R2794 VSS.n886 VSS.n885 75.4751
R2795 VSS.n889 VSS.n888 75.4751
R2796 VSS.n891 VSS.n890 75.4751
R2797 VSS.n894 VSS.n893 75.4751
R2798 VSS.n896 VSS.n895 75.4751
R2799 VSS.n899 VSS.n898 75.4751
R2800 VSS.n901 VSS.n900 75.4751
R2801 VSS.n904 VSS.n903 75.4751
R2802 VSS.n1885 VSS.n1535 75.2946
R2803 VSS.n1880 VSS.n1536 75.2946
R2804 VSS.n2110 VSS.n667 74.5417
R2805 VSS.n1640 VSS.n129 74.1652
R2806 VSS.n2019 VSS.n313 73.7435
R2807 VSS.t5 VSS.n2018 71.9877
R2808 VSS.n2027 VSS.t84 71.9877
R2809 VSS.n5 VSS.n3 70.8255
R2810 VSS.n83 VSS.n81 70.8255
R2811 VSS.n1090 VSS.n970 70.657
R2812 VSS.n907 VSS.n906 70.0483
R2813 VSS.n924 VSS.n923 70.0483
R2814 VSS.n917 VSS.n916 70.0483
R2815 VSS.n914 VSS.n913 70.0483
R2816 VSS.n1050 VSS.n1000 70.0401
R2817 VSS.n1006 VSS.n1004 70.0401
R2818 VSS.n1048 VSS.n1001 70.0054
R2819 VSS.n995 VSS.n993 70.0054
R2820 VSS.n1005 VSS.n1002 70.0054
R2821 VSS.n28 VSS.n27 69.6951
R2822 VSS.n85 VSS.n84 69.6951
R2823 VSS.n79 VSS.n78 69.6951
R2824 VSS.n1091 VSS.n968 69.6951
R2825 VSS.n1024 VSS.n1023 69.6951
R2826 VSS.n999 VSS.n996 69.6951
R2827 VSS.n1085 VSS.n1084 69.6951
R2828 VSS.n1089 VSS.n1088 69.6951
R2829 VSS.n5 VSS.n4 69.6895
R2830 VSS.n7 VSS.n6 69.6895
R2831 VSS.n50 VSS.n49 69.6895
R2832 VSS.n46 VSS.n45 69.6895
R2833 VSS.n39 VSS.n38 69.6895
R2834 VSS.n34 VSS.n33 69.6895
R2835 VSS.n95 VSS.n94 69.6895
R2836 VSS.n20 VSS.n19 69.6895
R2837 VSS.n105 VSS.n104 69.6895
R2838 VSS.n113 VSS.n112 69.6895
R2839 VSS.n116 VSS.n115 69.6895
R2840 VSS.n83 VSS.n82 69.6895
R2841 VSS.n44 VSS.n43 69.6895
R2842 VSS.n1093 VSS.n1092 69.6895
R2843 VSS.n1025 VSS.n1018 69.6895
R2844 VSS.n998 VSS.n997 69.6895
R2845 VSS.n992 VSS.n986 69.6895
R2846 VSS.n1083 VSS.n1082 69.6895
R2847 VSS.t89 VSS.n1522 68.4762
R2848 VSS.n461 VSS.t147 57.3715
R2849 VSS.n483 VSS.t186 57.3715
R2850 VSS.n525 VSS.n522 51.2005
R2851 VSS.n569 VSS.n566 51.2005
R2852 VSS.n1664 VSS.n1661 51.2005
R2853 VSS.n1708 VSS.n1705 51.2005
R2854 VSS.n1987 VSS.t89 50.9183
R2855 VSS.n1618 VSS.n9 48.7505
R2856 VSS.n1781 VSS.n1618 48.7505
R2857 VSS.n2019 VSS.t5 47.4067
R2858 VSS.t84 VSS.n2026 47.4067
R2859 VSS.n1506 VSS.n313 45.6509
R2860 VSS.n2336 VSS.n2335 45.2874
R2861 VSS.t64 VSS.n1526 43.8952
R2862 VSS.n2108 VSS.n2107 41.7429
R2863 VSS.n1496 VSS.n690 41.7429
R2864 VSS.t218 VSS.n1574 38.6169
R2865 VSS.n1830 VSS.t218 38.6169
R2866 VSS.n2226 VSS.n2225 36.1773
R2867 VSS.n1208 VSS.n671 36.1773
R2868 VSS.n1786 VSS.n1785 34.6377
R2869 VSS.n1776 VSS.n1774 34.6377
R2870 VSS.n1783 VSS.n1617 33.407
R2871 VSS.n1779 VSS.n1720 33.407
R2872 VSS.n1775 VSS.n1720 33.407
R2873 VSS.n1221 VSS.n812 30.1181
R2874 VSS.n1995 VSS.t3 26.3373
R2875 VSS.n1782 VSS.n1616 25.6631
R2876 VSS.n2382 VSS.n126 25.6631
R2877 VSS.n2376 VSS.n2375 25.6631
R2878 VSS.n2375 VSS.n2374 25.6631
R2879 VSS.n2374 VSS.n135 25.6631
R2880 VSS.n2368 VSS.n2367 25.6631
R2881 VSS.n2367 VSS.n2366 25.6631
R2882 VSS.n2360 VSS.n145 25.6631
R2883 VSS.n2360 VSS.n2359 25.6631
R2884 VSS.n2359 VSS.n2358 25.6631
R2885 VSS.n2352 VSS.n152 25.6631
R2886 VSS.n2352 VSS.n2351 25.6631
R2887 VSS.n2351 VSS.n2350 25.6631
R2888 VSS.n2344 VSS.n159 25.6631
R2889 VSS.n2344 VSS.n2343 25.6631
R2890 VSS.n2343 VSS.n2342 25.6631
R2891 VSS.n2336 VSS.n166 25.6631
R2892 VSS.n2223 VSS.n2222 25.6005
R2893 VSS.n2222 VSS.n2221 25.6005
R2894 VSS.n2221 VSS.n216 25.6005
R2895 VSS.n2215 VSS.n216 25.6005
R2896 VSS.n2215 VSS.n2214 25.6005
R2897 VSS.n2214 VSS.n2213 25.6005
R2898 VSS.n2213 VSS.n223 25.6005
R2899 VSS.n2207 VSS.n223 25.6005
R2900 VSS.n2207 VSS.n2206 25.6005
R2901 VSS.n2206 VSS.n2205 25.6005
R2902 VSS.n2205 VSS.n230 25.6005
R2903 VSS.n2199 VSS.n230 25.6005
R2904 VSS.n2199 VSS.n2198 25.6005
R2905 VSS.n2198 VSS.n2197 25.6005
R2906 VSS.n2197 VSS.n237 25.6005
R2907 VSS.n253 VSS.n237 25.6005
R2908 VSS.n254 VSS.n253 25.6005
R2909 VSS.n2184 VSS.n254 25.6005
R2910 VSS.n2184 VSS.n2183 25.6005
R2911 VSS.n2183 VSS.n2182 25.6005
R2912 VSS.n2182 VSS.n255 25.6005
R2913 VSS.n271 VSS.n255 25.6005
R2914 VSS.n2170 VSS.n271 25.6005
R2915 VSS.n2170 VSS.n2169 25.6005
R2916 VSS.n2169 VSS.n2168 25.6005
R2917 VSS.n2168 VSS.n272 25.6005
R2918 VSS.n287 VSS.n272 25.6005
R2919 VSS.n2156 VSS.n287 25.6005
R2920 VSS.n2156 VSS.n2155 25.6005
R2921 VSS.n2155 VSS.n2154 25.6005
R2922 VSS.n2154 VSS.n288 25.6005
R2923 VSS.n302 VSS.n288 25.6005
R2924 VSS.n2142 VSS.n302 25.6005
R2925 VSS.n2142 VSS.n2141 25.6005
R2926 VSS.n2141 VSS.n2140 25.6005
R2927 VSS.n2140 VSS.n303 25.6005
R2928 VSS.n318 VSS.n303 25.6005
R2929 VSS.n2128 VSS.n318 25.6005
R2930 VSS.n502 VSS.n215 25.6005
R2931 VSS.n505 VSS.n502 25.6005
R2932 VSS.n506 VSS.n505 25.6005
R2933 VSS.n509 VSS.n506 25.6005
R2934 VSS.n510 VSS.n509 25.6005
R2935 VSS.n513 VSS.n510 25.6005
R2936 VSS.n514 VSS.n513 25.6005
R2937 VSS.n517 VSS.n514 25.6005
R2938 VSS.n518 VSS.n517 25.6005
R2939 VSS.n521 VSS.n518 25.6005
R2940 VSS.n522 VSS.n521 25.6005
R2941 VSS.n526 VSS.n525 25.6005
R2942 VSS.n529 VSS.n526 25.6005
R2943 VSS.n530 VSS.n529 25.6005
R2944 VSS.n533 VSS.n530 25.6005
R2945 VSS.n534 VSS.n533 25.6005
R2946 VSS.n537 VSS.n534 25.6005
R2947 VSS.n538 VSS.n537 25.6005
R2948 VSS.n541 VSS.n538 25.6005
R2949 VSS.n542 VSS.n541 25.6005
R2950 VSS.n545 VSS.n542 25.6005
R2951 VSS.n546 VSS.n545 25.6005
R2952 VSS.n549 VSS.n546 25.6005
R2953 VSS.n550 VSS.n549 25.6005
R2954 VSS.n553 VSS.n550 25.6005
R2955 VSS.n554 VSS.n553 25.6005
R2956 VSS.n557 VSS.n554 25.6005
R2957 VSS.n558 VSS.n557 25.6005
R2958 VSS.n561 VSS.n558 25.6005
R2959 VSS.n562 VSS.n561 25.6005
R2960 VSS.n565 VSS.n562 25.6005
R2961 VSS.n566 VSS.n565 25.6005
R2962 VSS.n570 VSS.n569 25.6005
R2963 VSS.n573 VSS.n570 25.6005
R2964 VSS.n574 VSS.n573 25.6005
R2965 VSS.n577 VSS.n574 25.6005
R2966 VSS.n578 VSS.n577 25.6005
R2967 VSS.n581 VSS.n578 25.6005
R2968 VSS.n582 VSS.n581 25.6005
R2969 VSS.n585 VSS.n582 25.6005
R2970 VSS.n586 VSS.n585 25.6005
R2971 VSS.n591 VSS.n589 25.6005
R2972 VSS.n594 VSS.n592 25.6005
R2973 VSS.n595 VSS.n594 25.6005
R2974 VSS.n596 VSS.n595 25.6005
R2975 VSS.n597 VSS.n596 25.6005
R2976 VSS.n599 VSS.n597 25.6005
R2977 VSS.n600 VSS.n599 25.6005
R2978 VSS.n601 VSS.n600 25.6005
R2979 VSS.n602 VSS.n601 25.6005
R2980 VSS.n604 VSS.n602 25.6005
R2981 VSS.n605 VSS.n604 25.6005
R2982 VSS.n606 VSS.n605 25.6005
R2983 VSS.n607 VSS.n606 25.6005
R2984 VSS.n609 VSS.n607 25.6005
R2985 VSS.n610 VSS.n609 25.6005
R2986 VSS.n611 VSS.n610 25.6005
R2987 VSS.n612 VSS.n611 25.6005
R2988 VSS.n617 VSS.n612 25.6005
R2989 VSS.n618 VSS.n617 25.6005
R2990 VSS.n621 VSS.n618 25.6005
R2991 VSS.n622 VSS.n621 25.6005
R2992 VSS.n623 VSS.n622 25.6005
R2993 VSS.n626 VSS.n623 25.6005
R2994 VSS.n627 VSS.n626 25.6005
R2995 VSS.n630 VSS.n627 25.6005
R2996 VSS.n631 VSS.n630 25.6005
R2997 VSS.n632 VSS.n631 25.6005
R2998 VSS.n635 VSS.n632 25.6005
R2999 VSS.n636 VSS.n635 25.6005
R3000 VSS.n640 VSS.n636 25.6005
R3001 VSS.n641 VSS.n640 25.6005
R3002 VSS.n642 VSS.n641 25.6005
R3003 VSS.n647 VSS.n642 25.6005
R3004 VSS.n648 VSS.n647 25.6005
R3005 VSS.n651 VSS.n648 25.6005
R3006 VSS.n652 VSS.n651 25.6005
R3007 VSS.n653 VSS.n652 25.6005
R3008 VSS.n658 VSS.n653 25.6005
R3009 VSS.n659 VSS.n658 25.6005
R3010 VSS.n2127 VSS.n2126 25.6005
R3011 VSS.n2126 VSS.n319 25.6005
R3012 VSS.n345 VSS.n319 25.6005
R3013 VSS.n346 VSS.n345 25.6005
R3014 VSS.n349 VSS.n346 25.6005
R3015 VSS.n350 VSS.n349 25.6005
R3016 VSS.n353 VSS.n350 25.6005
R3017 VSS.n354 VSS.n353 25.6005
R3018 VSS.n357 VSS.n354 25.6005
R3019 VSS.n358 VSS.n357 25.6005
R3020 VSS.n361 VSS.n358 25.6005
R3021 VSS.n362 VSS.n361 25.6005
R3022 VSS.n365 VSS.n362 25.6005
R3023 VSS.n366 VSS.n365 25.6005
R3024 VSS.n369 VSS.n366 25.6005
R3025 VSS.n370 VSS.n369 25.6005
R3026 VSS.n373 VSS.n370 25.6005
R3027 VSS.n374 VSS.n373 25.6005
R3028 VSS.n377 VSS.n374 25.6005
R3029 VSS.n378 VSS.n377 25.6005
R3030 VSS.n381 VSS.n378 25.6005
R3031 VSS.n382 VSS.n381 25.6005
R3032 VSS.n385 VSS.n382 25.6005
R3033 VSS.n386 VSS.n385 25.6005
R3034 VSS.n389 VSS.n386 25.6005
R3035 VSS.n390 VSS.n389 25.6005
R3036 VSS.n393 VSS.n390 25.6005
R3037 VSS.n394 VSS.n393 25.6005
R3038 VSS.n397 VSS.n394 25.6005
R3039 VSS.n398 VSS.n397 25.6005
R3040 VSS.n401 VSS.n398 25.6005
R3041 VSS.n402 VSS.n401 25.6005
R3042 VSS.n405 VSS.n402 25.6005
R3043 VSS.n406 VSS.n405 25.6005
R3044 VSS.n409 VSS.n406 25.6005
R3045 VSS.n410 VSS.n409 25.6005
R3046 VSS.n413 VSS.n410 25.6005
R3047 VSS.n414 VSS.n413 25.6005
R3048 VSS.n417 VSS.n414 25.6005
R3049 VSS.n418 VSS.n417 25.6005
R3050 VSS.n421 VSS.n418 25.6005
R3051 VSS.n422 VSS.n421 25.6005
R3052 VSS.n425 VSS.n422 25.6005
R3053 VSS.n426 VSS.n425 25.6005
R3054 VSS.n429 VSS.n426 25.6005
R3055 VSS.n430 VSS.n429 25.6005
R3056 VSS.n660 VSS.n430 25.6005
R3057 VSS.n1981 VSS.n1528 25.6005
R3058 VSS.n1982 VSS.n1981 25.6005
R3059 VSS.n1983 VSS.n1982 25.6005
R3060 VSS.n1983 VSS.n1524 25.6005
R3061 VSS.n1989 VSS.n1524 25.6005
R3062 VSS.n1990 VSS.n1989 25.6005
R3063 VSS.n1991 VSS.n1990 25.6005
R3064 VSS.n1991 VSS.n1520 25.6005
R3065 VSS.n1997 VSS.n1520 25.6005
R3066 VSS.n1998 VSS.n1997 25.6005
R3067 VSS.n1999 VSS.n1998 25.6005
R3068 VSS.n1999 VSS.n1516 25.6005
R3069 VSS.n2005 VSS.n1516 25.6005
R3070 VSS.n2006 VSS.n2005 25.6005
R3071 VSS.n2007 VSS.n2006 25.6005
R3072 VSS.n2007 VSS.n1512 25.6005
R3073 VSS.n2013 VSS.n1512 25.6005
R3074 VSS.n2014 VSS.n2013 25.6005
R3075 VSS.n2015 VSS.n2014 25.6005
R3076 VSS.n2015 VSS.n1508 25.6005
R3077 VSS.n2021 VSS.n1508 25.6005
R3078 VSS.n2022 VSS.n2021 25.6005
R3079 VSS.n2023 VSS.n2022 25.6005
R3080 VSS.n2023 VSS.n1504 25.6005
R3081 VSS.n2029 VSS.n1504 25.6005
R3082 VSS.n2030 VSS.n2029 25.6005
R3083 VSS.n2031 VSS.n2030 25.6005
R3084 VSS.n2031 VSS.n1500 25.6005
R3085 VSS.n2037 VSS.n1500 25.6005
R3086 VSS.n2038 VSS.n2037 25.6005
R3087 VSS.n1907 VSS.n1906 25.6005
R3088 VSS.n1910 VSS.n1907 25.6005
R3089 VSS.n1911 VSS.n1910 25.6005
R3090 VSS.n1914 VSS.n1911 25.6005
R3091 VSS.n1915 VSS.n1914 25.6005
R3092 VSS.n1918 VSS.n1915 25.6005
R3093 VSS.n1919 VSS.n1918 25.6005
R3094 VSS.n1922 VSS.n1919 25.6005
R3095 VSS.n1923 VSS.n1922 25.6005
R3096 VSS.n1926 VSS.n1923 25.6005
R3097 VSS.n1927 VSS.n1926 25.6005
R3098 VSS.n1930 VSS.n1927 25.6005
R3099 VSS.n1931 VSS.n1930 25.6005
R3100 VSS.n1934 VSS.n1931 25.6005
R3101 VSS.n1935 VSS.n1934 25.6005
R3102 VSS.n1938 VSS.n1935 25.6005
R3103 VSS.n1939 VSS.n1938 25.6005
R3104 VSS.n1942 VSS.n1939 25.6005
R3105 VSS.n1943 VSS.n1942 25.6005
R3106 VSS.n1946 VSS.n1943 25.6005
R3107 VSS.n1947 VSS.n1946 25.6005
R3108 VSS.n1950 VSS.n1947 25.6005
R3109 VSS.n1951 VSS.n1950 25.6005
R3110 VSS.n1954 VSS.n1951 25.6005
R3111 VSS.n1955 VSS.n1954 25.6005
R3112 VSS.n1958 VSS.n1955 25.6005
R3113 VSS.n1960 VSS.n1958 25.6005
R3114 VSS.n1961 VSS.n1960 25.6005
R3115 VSS.n1974 VSS.n1961 25.6005
R3116 VSS.n1974 VSS.n1973 25.6005
R3117 VSS.n1973 VSS.n1972 25.6005
R3118 VSS.n1972 VSS.n1962 25.6005
R3119 VSS.n1967 VSS.n1962 25.6005
R3120 VSS.n1967 VSS.n1966 25.6005
R3121 VSS.n1966 VSS.n245 25.6005
R3122 VSS.n2191 VSS.n2190 25.6005
R3123 VSS.n2190 VSS.n2189 25.6005
R3124 VSS.n2189 VSS.n246 25.6005
R3125 VSS.n262 VSS.n246 25.6005
R3126 VSS.n2177 VSS.n262 25.6005
R3127 VSS.n2177 VSS.n2176 25.6005
R3128 VSS.n2176 VSS.n2175 25.6005
R3129 VSS.n2175 VSS.n263 25.6005
R3130 VSS.n279 VSS.n263 25.6005
R3131 VSS.n2163 VSS.n279 25.6005
R3132 VSS.n2163 VSS.n2162 25.6005
R3133 VSS.n2162 VSS.n2161 25.6005
R3134 VSS.n2161 VSS.n280 25.6005
R3135 VSS.n295 VSS.n280 25.6005
R3136 VSS.n2149 VSS.n295 25.6005
R3137 VSS.n2149 VSS.n2148 25.6005
R3138 VSS.n2148 VSS.n2147 25.6005
R3139 VSS.n2147 VSS.n296 25.6005
R3140 VSS.n310 VSS.n296 25.6005
R3141 VSS.n2135 VSS.n310 25.6005
R3142 VSS.n2135 VSS.n2134 25.6005
R3143 VSS.n2134 VSS.n2133 25.6005
R3144 VSS.n2133 VSS.n311 25.6005
R3145 VSS.n2120 VSS.n311 25.6005
R3146 VSS.n2120 VSS.n2119 25.6005
R3147 VSS.n2119 VSS.n2118 25.6005
R3148 VSS.n2118 VSS.n663 25.6005
R3149 VSS.n2112 VSS.n663 25.6005
R3150 VSS.n2112 VSS.n2111 25.6005
R3151 VSS.n2111 VSS.n2110 25.6005
R3152 VSS.n2089 VSS.n2088 25.6005
R3153 VSS.n2088 VSS.n2087 25.6005
R3154 VSS.n2087 VSS.n2086 25.6005
R3155 VSS.n2086 VSS.n2084 25.6005
R3156 VSS.n2084 VSS.n2081 25.6005
R3157 VSS.n2081 VSS.n2080 25.6005
R3158 VSS.n2080 VSS.n2077 25.6005
R3159 VSS.n2077 VSS.n2076 25.6005
R3160 VSS.n2076 VSS.n2073 25.6005
R3161 VSS.n2073 VSS.n2072 25.6005
R3162 VSS.n2072 VSS.n2069 25.6005
R3163 VSS.n2069 VSS.n2068 25.6005
R3164 VSS.n2068 VSS.n2065 25.6005
R3165 VSS.n2065 VSS.n2064 25.6005
R3166 VSS.n2064 VSS.n2061 25.6005
R3167 VSS.n2061 VSS.n2060 25.6005
R3168 VSS.n2060 VSS.n2057 25.6005
R3169 VSS.n2057 VSS.n2056 25.6005
R3170 VSS.n2056 VSS.n2053 25.6005
R3171 VSS.n2053 VSS.n2052 25.6005
R3172 VSS.n2052 VSS.n2049 25.6005
R3173 VSS.n2049 VSS.n2048 25.6005
R3174 VSS.n2048 VSS.n2045 25.6005
R3175 VSS.n2045 VSS.n2044 25.6005
R3176 VSS.n2044 VSS.n2041 25.6005
R3177 VSS.n2041 VSS.n2040 25.6005
R3178 VSS.n2040 VSS.n675 25.6005
R3179 VSS.n2095 VSS.n675 25.6005
R3180 VSS.n2096 VSS.n2095 25.6005
R3181 VSS.n2104 VSS.n2096 25.6005
R3182 VSS.n2104 VSS.n2103 25.6005
R3183 VSS.n2103 VSS.n2102 25.6005
R3184 VSS.n2102 VSS.n2101 25.6005
R3185 VSS.n2101 VSS.n2099 25.6005
R3186 VSS.n2099 VSS.n2097 25.6005
R3187 VSS.n1874 VSS.n1535 25.6005
R3188 VSS.n1874 VSS.n1873 25.6005
R3189 VSS.n1873 VSS.n1872 25.6005
R3190 VSS.n1872 VSS.n1541 25.6005
R3191 VSS.n1866 VSS.n1541 25.6005
R3192 VSS.n1866 VSS.n1865 25.6005
R3193 VSS.n1865 VSS.n1864 25.6005
R3194 VSS.n1864 VSS.n1548 25.6005
R3195 VSS.n1858 VSS.n1548 25.6005
R3196 VSS.n1858 VSS.n1857 25.6005
R3197 VSS.n1857 VSS.n1856 25.6005
R3198 VSS.n1856 VSS.n1555 25.6005
R3199 VSS.n1850 VSS.n1555 25.6005
R3200 VSS.n1850 VSS.n1849 25.6005
R3201 VSS.n1849 VSS.n1848 25.6005
R3202 VSS.n1848 VSS.n1562 25.6005
R3203 VSS.n1842 VSS.n1562 25.6005
R3204 VSS.n1842 VSS.n1841 25.6005
R3205 VSS.n1841 VSS.n1840 25.6005
R3206 VSS.n1840 VSS.n1569 25.6005
R3207 VSS.n1834 VSS.n1569 25.6005
R3208 VSS.n1834 VSS.n1833 25.6005
R3209 VSS.n1833 VSS.n1832 25.6005
R3210 VSS.n1832 VSS.n1576 25.6005
R3211 VSS.n1826 VSS.n1576 25.6005
R3212 VSS.n1826 VSS.n1825 25.6005
R3213 VSS.n1825 VSS.n1824 25.6005
R3214 VSS.n1824 VSS.n1583 25.6005
R3215 VSS.n1818 VSS.n1583 25.6005
R3216 VSS.n1818 VSS.n1817 25.6005
R3217 VSS.n1817 VSS.n1816 25.6005
R3218 VSS.n1816 VSS.n1590 25.6005
R3219 VSS.n1810 VSS.n1590 25.6005
R3220 VSS.n1810 VSS.n1809 25.6005
R3221 VSS.n1809 VSS.n1808 25.6005
R3222 VSS.n1808 VSS.n1597 25.6005
R3223 VSS.n1802 VSS.n1597 25.6005
R3224 VSS.n1802 VSS.n1801 25.6005
R3225 VSS.n1801 VSS.n1800 25.6005
R3226 VSS.n1800 VSS.n1604 25.6005
R3227 VSS.n1794 VSS.n1604 25.6005
R3228 VSS.n1794 VSS.n1793 25.6005
R3229 VSS.n1793 VSS.n1792 25.6005
R3230 VSS.n1792 VSS.n1611 25.6005
R3231 VSS.n1786 VSS.n1611 25.6005
R3232 VSS.n1885 VSS.n1884 25.6005
R3233 VSS.n1884 VSS.n1883 25.6005
R3234 VSS.n1883 VSS.n1882 25.6005
R3235 VSS.n1882 VSS.n1880 25.6005
R3236 VSS.n1538 VSS.n1536 25.6005
R3237 VSS.n1721 VSS.n1538 25.6005
R3238 VSS.n1722 VSS.n1721 25.6005
R3239 VSS.n1723 VSS.n1722 25.6005
R3240 VSS.n1724 VSS.n1723 25.6005
R3241 VSS.n1726 VSS.n1724 25.6005
R3242 VSS.n1727 VSS.n1726 25.6005
R3243 VSS.n1728 VSS.n1727 25.6005
R3244 VSS.n1729 VSS.n1728 25.6005
R3245 VSS.n1731 VSS.n1729 25.6005
R3246 VSS.n1732 VSS.n1731 25.6005
R3247 VSS.n1733 VSS.n1732 25.6005
R3248 VSS.n1734 VSS.n1733 25.6005
R3249 VSS.n1736 VSS.n1734 25.6005
R3250 VSS.n1737 VSS.n1736 25.6005
R3251 VSS.n1738 VSS.n1737 25.6005
R3252 VSS.n1739 VSS.n1738 25.6005
R3253 VSS.n1741 VSS.n1739 25.6005
R3254 VSS.n1742 VSS.n1741 25.6005
R3255 VSS.n1743 VSS.n1742 25.6005
R3256 VSS.n1744 VSS.n1743 25.6005
R3257 VSS.n1746 VSS.n1744 25.6005
R3258 VSS.n1747 VSS.n1746 25.6005
R3259 VSS.n1748 VSS.n1747 25.6005
R3260 VSS.n1749 VSS.n1748 25.6005
R3261 VSS.n1751 VSS.n1749 25.6005
R3262 VSS.n1752 VSS.n1751 25.6005
R3263 VSS.n1753 VSS.n1752 25.6005
R3264 VSS.n1754 VSS.n1753 25.6005
R3265 VSS.n1756 VSS.n1754 25.6005
R3266 VSS.n1757 VSS.n1756 25.6005
R3267 VSS.n1758 VSS.n1757 25.6005
R3268 VSS.n1759 VSS.n1758 25.6005
R3269 VSS.n1761 VSS.n1759 25.6005
R3270 VSS.n1762 VSS.n1761 25.6005
R3271 VSS.n1763 VSS.n1762 25.6005
R3272 VSS.n1764 VSS.n1763 25.6005
R3273 VSS.n1766 VSS.n1764 25.6005
R3274 VSS.n1767 VSS.n1766 25.6005
R3275 VSS.n1768 VSS.n1767 25.6005
R3276 VSS.n1769 VSS.n1768 25.6005
R3277 VSS.n1771 VSS.n1769 25.6005
R3278 VSS.n1772 VSS.n1771 25.6005
R3279 VSS.n1773 VSS.n1772 25.6005
R3280 VSS.n1774 VSS.n1773 25.6005
R3281 VSS.n2380 VSS.n129 25.6005
R3282 VSS.n2380 VSS.n2379 25.6005
R3283 VSS.n2379 VSS.n2378 25.6005
R3284 VSS.n2378 VSS.n130 25.6005
R3285 VSS.n2372 VSS.n130 25.6005
R3286 VSS.n2372 VSS.n2371 25.6005
R3287 VSS.n2371 VSS.n2370 25.6005
R3288 VSS.n2370 VSS.n137 25.6005
R3289 VSS.n2364 VSS.n137 25.6005
R3290 VSS.n2364 VSS.n2363 25.6005
R3291 VSS.n2363 VSS.n2362 25.6005
R3292 VSS.n2362 VSS.n143 25.6005
R3293 VSS.n2356 VSS.n143 25.6005
R3294 VSS.n2356 VSS.n2355 25.6005
R3295 VSS.n2355 VSS.n2354 25.6005
R3296 VSS.n2354 VSS.n150 25.6005
R3297 VSS.n2348 VSS.n150 25.6005
R3298 VSS.n2348 VSS.n2347 25.6005
R3299 VSS.n2347 VSS.n2346 25.6005
R3300 VSS.n2346 VSS.n157 25.6005
R3301 VSS.n2340 VSS.n157 25.6005
R3302 VSS.n2340 VSS.n2339 25.6005
R3303 VSS.n2339 VSS.n2338 25.6005
R3304 VSS.n1641 VSS.n1640 25.6005
R3305 VSS.n1644 VSS.n1641 25.6005
R3306 VSS.n1645 VSS.n1644 25.6005
R3307 VSS.n1648 VSS.n1645 25.6005
R3308 VSS.n1649 VSS.n1648 25.6005
R3309 VSS.n1652 VSS.n1649 25.6005
R3310 VSS.n1653 VSS.n1652 25.6005
R3311 VSS.n1656 VSS.n1653 25.6005
R3312 VSS.n1657 VSS.n1656 25.6005
R3313 VSS.n1660 VSS.n1657 25.6005
R3314 VSS.n1661 VSS.n1660 25.6005
R3315 VSS.n1665 VSS.n1664 25.6005
R3316 VSS.n1668 VSS.n1665 25.6005
R3317 VSS.n1669 VSS.n1668 25.6005
R3318 VSS.n1672 VSS.n1669 25.6005
R3319 VSS.n1673 VSS.n1672 25.6005
R3320 VSS.n1676 VSS.n1673 25.6005
R3321 VSS.n1677 VSS.n1676 25.6005
R3322 VSS.n1680 VSS.n1677 25.6005
R3323 VSS.n1681 VSS.n1680 25.6005
R3324 VSS.n1684 VSS.n1681 25.6005
R3325 VSS.n1685 VSS.n1684 25.6005
R3326 VSS.n1688 VSS.n1685 25.6005
R3327 VSS.n1689 VSS.n1688 25.6005
R3328 VSS.n1692 VSS.n1689 25.6005
R3329 VSS.n1693 VSS.n1692 25.6005
R3330 VSS.n1696 VSS.n1693 25.6005
R3331 VSS.n1697 VSS.n1696 25.6005
R3332 VSS.n1700 VSS.n1697 25.6005
R3333 VSS.n1701 VSS.n1700 25.6005
R3334 VSS.n1704 VSS.n1701 25.6005
R3335 VSS.n1705 VSS.n1704 25.6005
R3336 VSS.n1709 VSS.n1708 25.6005
R3337 VSS.n1712 VSS.n1709 25.6005
R3338 VSS.n1713 VSS.n1712 25.6005
R3339 VSS.n1714 VSS.n1713 25.6005
R3340 VSS.n1714 VSS.n121 25.6005
R3341 VSS.n2384 VSS.n122 25.6005
R3342 VSS.n2228 VSS.n122 25.6005
R3343 VSS.n2229 VSS.n2228 25.6005
R3344 VSS.n2230 VSS.n2229 25.6005
R3345 VSS.n2232 VSS.n2230 25.6005
R3346 VSS.n2233 VSS.n2232 25.6005
R3347 VSS.n2234 VSS.n2233 25.6005
R3348 VSS.n2235 VSS.n2234 25.6005
R3349 VSS.n2237 VSS.n2235 25.6005
R3350 VSS.n2238 VSS.n2237 25.6005
R3351 VSS.n2239 VSS.n2238 25.6005
R3352 VSS.n2240 VSS.n2239 25.6005
R3353 VSS.n2242 VSS.n2240 25.6005
R3354 VSS.n2243 VSS.n2242 25.6005
R3355 VSS.n2244 VSS.n2243 25.6005
R3356 VSS.n2245 VSS.n2244 25.6005
R3357 VSS.n2247 VSS.n2245 25.6005
R3358 VSS.n2248 VSS.n2247 25.6005
R3359 VSS.n2249 VSS.n2248 25.6005
R3360 VSS.n2250 VSS.n2249 25.6005
R3361 VSS.n2252 VSS.n2250 25.6005
R3362 VSS.n2253 VSS.n2252 25.6005
R3363 VSS.n2332 VSS.n164 25.6005
R3364 VSS.n2332 VSS.n2331 25.6005
R3365 VSS.n2331 VSS.n2330 25.6005
R3366 VSS.n2330 VSS.n2328 25.6005
R3367 VSS.n2328 VSS.n2325 25.6005
R3368 VSS.n2325 VSS.n2324 25.6005
R3369 VSS.n2324 VSS.n2321 25.6005
R3370 VSS.n2321 VSS.n2320 25.6005
R3371 VSS.n2320 VSS.n2317 25.6005
R3372 VSS.n2317 VSS.n2316 25.6005
R3373 VSS.n2316 VSS.n2313 25.6005
R3374 VSS.n2313 VSS.n2312 25.6005
R3375 VSS.n2312 VSS.n2309 25.6005
R3376 VSS.n2309 VSS.n2308 25.6005
R3377 VSS.n2308 VSS.n2305 25.6005
R3378 VSS.n2305 VSS.n2304 25.6005
R3379 VSS.n2304 VSS.n2301 25.6005
R3380 VSS.n2301 VSS.n2300 25.6005
R3381 VSS.n2300 VSS.n2297 25.6005
R3382 VSS.n2297 VSS.n2296 25.6005
R3383 VSS.n2296 VSS.n2293 25.6005
R3384 VSS.n2293 VSS.n2292 25.6005
R3385 VSS.n2292 VSS.n2289 25.6005
R3386 VSS.n2289 VSS.n2288 25.6005
R3387 VSS.n2288 VSS.n2285 25.6005
R3388 VSS.n2285 VSS.n2284 25.6005
R3389 VSS.n2284 VSS.n2281 25.6005
R3390 VSS.n2281 VSS.n2280 25.6005
R3391 VSS.n2280 VSS.n2277 25.6005
R3392 VSS.n2277 VSS.n2276 25.6005
R3393 VSS.n2276 VSS.n2273 25.6005
R3394 VSS.n2273 VSS.n2272 25.6005
R3395 VSS.n2272 VSS.n2269 25.6005
R3396 VSS.n2269 VSS.n2268 25.6005
R3397 VSS.n2268 VSS.n2265 25.6005
R3398 VSS.n2265 VSS.n2264 25.6005
R3399 VSS.n2264 VSS.n2261 25.6005
R3400 VSS.n2261 VSS.n2260 25.6005
R3401 VSS.n2260 VSS.n2257 25.6005
R3402 VSS.n2257 VSS.n2256 25.6005
R3403 VSS.n2256 VSS.n2254 25.6005
R3404 VSS.n1206 VSS.n819 25.6005
R3405 VSS.n1219 VSS.n819 25.6005
R3406 VSS.n1220 VSS.n1219 25.6005
R3407 VSS.n1221 VSS.n1220 25.6005
R3408 VSS.n1233 VSS.n812 25.6005
R3409 VSS.n1234 VSS.n1233 25.6005
R3410 VSS.n1235 VSS.n1234 25.6005
R3411 VSS.n1235 VSS.n804 25.6005
R3412 VSS.n1245 VSS.n804 25.6005
R3413 VSS.n1246 VSS.n1245 25.6005
R3414 VSS.n1247 VSS.n1246 25.6005
R3415 VSS.n1247 VSS.n796 25.6005
R3416 VSS.n1257 VSS.n796 25.6005
R3417 VSS.n1258 VSS.n1257 25.6005
R3418 VSS.n1259 VSS.n1258 25.6005
R3419 VSS.n1259 VSS.n788 25.6005
R3420 VSS.n1269 VSS.n788 25.6005
R3421 VSS.n1270 VSS.n1269 25.6005
R3422 VSS.n1271 VSS.n1270 25.6005
R3423 VSS.n1271 VSS.n780 25.6005
R3424 VSS.n1281 VSS.n780 25.6005
R3425 VSS.n1282 VSS.n1281 25.6005
R3426 VSS.n1283 VSS.n1282 25.6005
R3427 VSS.n1283 VSS.n772 25.6005
R3428 VSS.n1293 VSS.n772 25.6005
R3429 VSS.n1294 VSS.n1293 25.6005
R3430 VSS.n1295 VSS.n1294 25.6005
R3431 VSS.n1295 VSS.n764 25.6005
R3432 VSS.n1305 VSS.n764 25.6005
R3433 VSS.n1306 VSS.n1305 25.6005
R3434 VSS.n1307 VSS.n1306 25.6005
R3435 VSS.n1307 VSS.n756 25.6005
R3436 VSS.n1317 VSS.n756 25.6005
R3437 VSS.n1318 VSS.n1317 25.6005
R3438 VSS.n1319 VSS.n1318 25.6005
R3439 VSS.n1319 VSS.n748 25.6005
R3440 VSS.n1330 VSS.n748 25.6005
R3441 VSS.n1331 VSS.n1330 25.6005
R3442 VSS.n1332 VSS.n1331 25.6005
R3443 VSS.n1332 VSS.n741 25.6005
R3444 VSS.n1343 VSS.n741 25.6005
R3445 VSS.n1344 VSS.n1343 25.6005
R3446 VSS.n1345 VSS.n1344 25.6005
R3447 VSS.n1345 VSS.n734 25.6005
R3448 VSS.n1356 VSS.n734 25.6005
R3449 VSS.n1357 VSS.n1356 25.6005
R3450 VSS.n1358 VSS.n1357 25.6005
R3451 VSS.n1358 VSS.n727 25.6005
R3452 VSS.n1370 VSS.n727 25.6005
R3453 VSS.n1371 VSS.n1370 25.6005
R3454 VSS.n1372 VSS.n1371 25.6005
R3455 VSS.n1372 VSS.n723 25.6005
R3456 VSS.n1493 VSS.n1492 25.6005
R3457 VSS.n1492 VSS.n1491 25.6005
R3458 VSS.n1491 VSS.n1490 25.6005
R3459 VSS.n1490 VSS.n1488 25.6005
R3460 VSS.n1488 VSS.n1485 25.6005
R3461 VSS.n1485 VSS.n1484 25.6005
R3462 VSS.n1484 VSS.n1481 25.6005
R3463 VSS.n1481 VSS.n1480 25.6005
R3464 VSS.n1480 VSS.n1477 25.6005
R3465 VSS.n1477 VSS.n1476 25.6005
R3466 VSS.n1476 VSS.n1473 25.6005
R3467 VSS.n1473 VSS.n1472 25.6005
R3468 VSS.n1472 VSS.n1469 25.6005
R3469 VSS.n1469 VSS.n1468 25.6005
R3470 VSS.n1468 VSS.n1465 25.6005
R3471 VSS.n1465 VSS.n1464 25.6005
R3472 VSS.n1464 VSS.n1461 25.6005
R3473 VSS.n1461 VSS.n1460 25.6005
R3474 VSS.n1460 VSS.n1457 25.6005
R3475 VSS.n1457 VSS.n1456 25.6005
R3476 VSS.n1456 VSS.n1453 25.6005
R3477 VSS.n1453 VSS.n1452 25.6005
R3478 VSS.n1452 VSS.n1449 25.6005
R3479 VSS.n1449 VSS.n1448 25.6005
R3480 VSS.n1448 VSS.n1445 25.6005
R3481 VSS.n1445 VSS.n1444 25.6005
R3482 VSS.n1444 VSS.n1441 25.6005
R3483 VSS.n1441 VSS.n1440 25.6005
R3484 VSS.n1440 VSS.n1437 25.6005
R3485 VSS.n1437 VSS.n1436 25.6005
R3486 VSS.n1436 VSS.n1433 25.6005
R3487 VSS.n1433 VSS.n1432 25.6005
R3488 VSS.n1432 VSS.n1429 25.6005
R3489 VSS.n1429 VSS.n1428 25.6005
R3490 VSS.n1428 VSS.n1425 25.6005
R3491 VSS.n1425 VSS.n1424 25.6005
R3492 VSS.n1424 VSS.n1421 25.6005
R3493 VSS.n1421 VSS.n1420 25.6005
R3494 VSS.n1420 VSS.n1417 25.6005
R3495 VSS.n1417 VSS.n1416 25.6005
R3496 VSS.n1416 VSS.n1413 25.6005
R3497 VSS.n1413 VSS.n1412 25.6005
R3498 VSS.n1412 VSS.n1409 25.6005
R3499 VSS.n1409 VSS.n1408 25.6005
R3500 VSS.n1408 VSS.n1405 25.6005
R3501 VSS.n1405 VSS.n1404 25.6005
R3502 VSS.n1404 VSS.n1401 25.6005
R3503 VSS.n1401 VSS.n1400 25.6005
R3504 VSS.n1400 VSS.n1397 25.6005
R3505 VSS.n1397 VSS.n1396 25.6005
R3506 VSS.n1396 VSS.n1393 25.6005
R3507 VSS.n1393 VSS.n1392 25.6005
R3508 VSS.n1392 VSS.n1389 25.6005
R3509 VSS.n1389 VSS.n1388 25.6005
R3510 VSS.n1388 VSS.n1385 25.6005
R3511 VSS.n1385 VSS.n1384 25.6005
R3512 VSS.n1384 VSS.n1381 25.6005
R3513 VSS.n1381 VSS.n1380 25.6005
R3514 VSS.n1380 VSS.n1378 25.6005
R3515 VSS.n1213 VSS.n1212 25.6005
R3516 VSS.n1214 VSS.n1213 25.6005
R3517 VSS.n1214 VSS.n815 25.6005
R3518 VSS.n1227 VSS.n815 25.6005
R3519 VSS.n1228 VSS.n1227 25.6005
R3520 VSS.n1229 VSS.n1228 25.6005
R3521 VSS.n1229 VSS.n807 25.6005
R3522 VSS.n1239 VSS.n807 25.6005
R3523 VSS.n1240 VSS.n1239 25.6005
R3524 VSS.n1241 VSS.n1240 25.6005
R3525 VSS.n1241 VSS.n799 25.6005
R3526 VSS.n1251 VSS.n799 25.6005
R3527 VSS.n1252 VSS.n1251 25.6005
R3528 VSS.n1253 VSS.n1252 25.6005
R3529 VSS.n1253 VSS.n791 25.6005
R3530 VSS.n1263 VSS.n791 25.6005
R3531 VSS.n1264 VSS.n1263 25.6005
R3532 VSS.n1265 VSS.n1264 25.6005
R3533 VSS.n1265 VSS.n784 25.6005
R3534 VSS.n1275 VSS.n784 25.6005
R3535 VSS.n1276 VSS.n1275 25.6005
R3536 VSS.n1277 VSS.n1276 25.6005
R3537 VSS.n1277 VSS.n776 25.6005
R3538 VSS.n1287 VSS.n776 25.6005
R3539 VSS.n1288 VSS.n1287 25.6005
R3540 VSS.n1289 VSS.n1288 25.6005
R3541 VSS.n1289 VSS.n768 25.6005
R3542 VSS.n1299 VSS.n768 25.6005
R3543 VSS.n1300 VSS.n1299 25.6005
R3544 VSS.n1301 VSS.n1300 25.6005
R3545 VSS.n1301 VSS.n760 25.6005
R3546 VSS.n1311 VSS.n760 25.6005
R3547 VSS.n1312 VSS.n1311 25.6005
R3548 VSS.n1313 VSS.n1312 25.6005
R3549 VSS.n1313 VSS.n752 25.6005
R3550 VSS.n1323 VSS.n752 25.6005
R3551 VSS.n1324 VSS.n1323 25.6005
R3552 VSS.n1325 VSS.n1324 25.6005
R3553 VSS.n1325 VSS.n745 25.6005
R3554 VSS.n1336 VSS.n745 25.6005
R3555 VSS.n1337 VSS.n1336 25.6005
R3556 VSS.n1338 VSS.n1337 25.6005
R3557 VSS.n1338 VSS.n738 25.6005
R3558 VSS.n1349 VSS.n738 25.6005
R3559 VSS.n1350 VSS.n1349 25.6005
R3560 VSS.n1351 VSS.n1350 25.6005
R3561 VSS.n1351 VSS.n731 25.6005
R3562 VSS.n1362 VSS.n731 25.6005
R3563 VSS.n1363 VSS.n1362 25.6005
R3564 VSS.n1365 VSS.n1363 25.6005
R3565 VSS.n1365 VSS.n1364 25.6005
R3566 VSS.n1364 VSS.n724 25.6005
R3567 VSS.n1377 VSS.n724 25.6005
R3568 VSS.n1205 VSS.n1204 25.6005
R3569 VSS.n1204 VSS.n827 25.6005
R3570 VSS.n1199 VSS.n827 25.6005
R3571 VSS.n1199 VSS.n1198 25.6005
R3572 VSS.n1198 VSS.n1197 25.6005
R3573 VSS.n1197 VSS.n830 25.6005
R3574 VSS.n1192 VSS.n830 25.6005
R3575 VSS.n1192 VSS.n1191 25.6005
R3576 VSS.n1191 VSS.n1190 25.6005
R3577 VSS.n1190 VSS.n833 25.6005
R3578 VSS.n1185 VSS.n833 25.6005
R3579 VSS.n1185 VSS.n1184 25.6005
R3580 VSS.n1184 VSS.n1183 25.6005
R3581 VSS.n1183 VSS.n836 25.6005
R3582 VSS.n1178 VSS.n836 25.6005
R3583 VSS.n1178 VSS.n1177 25.6005
R3584 VSS.n1177 VSS.n1176 25.6005
R3585 VSS.n1176 VSS.n839 25.6005
R3586 VSS.n1171 VSS.n839 25.6005
R3587 VSS.n1171 VSS.n1170 25.6005
R3588 VSS.n1170 VSS.n1169 25.6005
R3589 VSS.n1169 VSS.n842 25.6005
R3590 VSS.n1164 VSS.n842 25.6005
R3591 VSS.n1164 VSS.n1163 25.6005
R3592 VSS.n1163 VSS.n1162 25.6005
R3593 VSS.n1162 VSS.n845 25.6005
R3594 VSS.n1157 VSS.n845 25.6005
R3595 VSS.n1157 VSS.n1156 25.6005
R3596 VSS.n1156 VSS.n1155 25.6005
R3597 VSS.n1155 VSS.n848 25.6005
R3598 VSS.n1150 VSS.n848 25.6005
R3599 VSS.n1150 VSS.n1149 25.6005
R3600 VSS.n1149 VSS.n1148 25.6005
R3601 VSS.n1148 VSS.n851 25.6005
R3602 VSS.n1143 VSS.n851 25.6005
R3603 VSS.n1143 VSS.n1142 25.6005
R3604 VSS.n1142 VSS.n1141 25.6005
R3605 VSS.n1141 VSS.n854 25.6005
R3606 VSS.n1136 VSS.n854 25.6005
R3607 VSS.n1136 VSS.n1135 25.6005
R3608 VSS.n1135 VSS.n1134 25.6005
R3609 VSS.n1134 VSS.n857 25.6005
R3610 VSS.n1129 VSS.n857 25.6005
R3611 VSS.n1129 VSS.n1128 25.6005
R3612 VSS.n1128 VSS.n1127 25.6005
R3613 VSS.n1127 VSS.n860 25.6005
R3614 VSS.n1122 VSS.n860 25.6005
R3615 VSS.n1122 VSS.n1121 25.6005
R3616 VSS.n1121 VSS.n1120 25.6005
R3617 VSS.n1120 VSS.n863 25.6005
R3618 VSS.n1115 VSS.n863 25.6005
R3619 VSS.n1115 VSS.n1114 25.6005
R3620 VSS.n1114 VSS.n1113 25.6005
R3621 VSS.n1113 VSS.n866 25.6005
R3622 VSS.n1108 VSS.n866 25.6005
R3623 VSS.n1108 VSS.n1107 25.6005
R3624 VSS.n1107 VSS.n1106 25.6005
R3625 VSS.n1106 VSS.n1101 25.6005
R3626 VSS.n2368 VSS.t216 25.2857
R3627 VSS.n1779 VSS.n1618 25.0554
R3628 VSS.n586 VSS.n501 24.4711
R3629 VSS.n2225 VSS.n212 23.6545
R3630 VSS.n2219 VSS.n212 23.6545
R3631 VSS.n2218 VSS.n2217 23.6545
R3632 VSS.n2217 VSS.n221 23.6545
R3633 VSS.n2211 VSS.n2210 23.6545
R3634 VSS.n2210 VSS.n2209 23.6545
R3635 VSS.n2209 VSS.n228 23.6545
R3636 VSS.n2203 VSS.n2202 23.6545
R3637 VSS.n2202 VSS.n2201 23.6545
R3638 VSS.n2201 VSS.n235 23.6545
R3639 VSS.n2195 VSS.n2194 23.6545
R3640 VSS.n2116 VSS.n665 23.6545
R3641 VSS.n2116 VSS.n2115 23.6545
R3642 VSS.n2115 VSS.n2114 23.6545
R3643 VSS.n2108 VSS.n669 23.6545
R3644 VSS.n1225 VSS.n1224 23.6545
R3645 VSS.n1231 VSS.n809 23.6545
R3646 VSS.n1237 VSS.n809 23.6545
R3647 VSS.n1237 VSS.n810 23.6545
R3648 VSS.n1243 VSS.n801 23.6545
R3649 VSS.n1249 VSS.n801 23.6545
R3650 VSS.n1249 VSS.n802 23.6545
R3651 VSS.n1255 VSS.n793 23.6545
R3652 VSS.n1261 VSS.n793 23.6545
R3653 VSS.n1261 VSS.n794 23.6545
R3654 VSS.n1267 VSS.n786 23.6545
R3655 VSS.n1273 VSS.n786 23.6545
R3656 VSS.n1279 VSS.n782 23.6545
R3657 VSS.n1279 VSS.n778 23.6545
R3658 VSS.n1285 VSS.n778 23.6545
R3659 VSS.n1291 VSS.n774 23.6545
R3660 VSS.n1291 VSS.n770 23.6545
R3661 VSS.n1297 VSS.n770 23.6545
R3662 VSS.n1303 VSS.n766 23.6545
R3663 VSS.n1303 VSS.n762 23.6545
R3664 VSS.n1309 VSS.n762 23.6545
R3665 VSS.n1315 VSS.n758 23.6545
R3666 VSS.n1315 VSS.n754 23.6545
R3667 VSS.n1321 VSS.n754 23.6545
R3668 VSS.n1328 VSS.n750 23.6545
R3669 VSS.n1328 VSS.n1327 23.6545
R3670 VSS.n1334 VSS.n743 23.6545
R3671 VSS.n1341 VSS.n743 23.6545
R3672 VSS.n1341 VSS.n1340 23.6545
R3673 VSS.n1347 VSS.n736 23.6545
R3674 VSS.n1354 VSS.n736 23.6545
R3675 VSS.n1354 VSS.n1353 23.6545
R3676 VSS.n1360 VSS.n729 23.6545
R3677 VSS.n1368 VSS.n729 23.6545
R3678 VSS.n1368 VSS.n1367 23.6545
R3679 VSS.n1374 VSS.n690 23.6545
R3680 VSS.t20 VSS.n750 23.3067
R3681 VSS.n2011 VSS.t2 22.8257
R3682 VSS.t61 VSS.n2034 22.8257
R3683 VSS.t27 VSS.n2218 22.611
R3684 VSS.n1267 VSS.t17 22.611
R3685 VSS.n2194 VSS.n2193 21.9153
R3686 VSS.n614 VSS.n242 21.9153
R3687 VSS.n2186 VSS.n249 21.9153
R3688 VSS.n619 VSS.n257 21.9153
R3689 VSS.n2180 VSS.n2179 21.9153
R3690 VSS.n2173 VSS.n266 21.9153
R3691 VSS.n2172 VSS.n268 21.9153
R3692 VSS.n282 VSS.n276 21.9153
R3693 VSS.n2159 VSS.n283 21.9153
R3694 VSS.n638 VSS.n290 21.9153
R3695 VSS.n2152 VSS.n2151 21.9153
R3696 VSS.n644 VSS.n292 21.9153
R3697 VSS.n2144 VSS.n299 21.9153
R3698 VSS.n649 VSS.n305 21.9153
R3699 VSS.n2138 VSS.n2137 21.9153
R3700 VSS.n2130 VSS.n315 21.9153
R3701 VSS.n1719 VSS.n1717 20.757
R3702 VSS.n2366 VSS.t215 20.757
R3703 VSS.n166 VSS.t30 20.757
R3704 VSS.n2376 VSS.t22 20.0022
R3705 VSS.t10 VSS.n221 19.8282
R3706 VSS.n2123 VSS.n315 19.8282
R3707 VSS.n1273 VSS.t6 19.8282
R3708 VSS.n1210 VSS.n1209 19.4803
R3709 VSS.n1217 VSS.n821 19.4803
R3710 VSS.n1216 VSS.n822 19.4803
R3711 VSS.n1223 VSS.n817 19.4803
R3712 VSS.n1781 VSS.n1780 19.2474
R3713 VSS.n1100 VSS.n824 19.2005
R3714 VSS.n628 VSS.t1 19.1324
R3715 VSS.n669 VSS.t102 19.1324
R3716 VSS.n1327 VSS.t12 19.1324
R3717 VSS.n1374 VSS.t38 19.1324
R3718 VSS.t313 VSS.n2165 18.4367
R3719 VSS.t19 VSS.n758 18.4367
R3720 VSS.n1255 VSS.t15 17.741
R3721 VSS.n431 VSS.t278 17.4005
R3722 VSS.n431 VSS.t273 17.4005
R3723 VSS.n432 VSS.t235 17.4005
R3724 VSS.n432 VSS.t229 17.4005
R3725 VSS.n434 VSS.t222 17.4005
R3726 VSS.n434 VSS.t274 17.4005
R3727 VSS.n435 VSS.t297 17.4005
R3728 VSS.n435 VSS.t234 17.4005
R3729 VSS.n438 VSS.t275 17.4005
R3730 VSS.n438 VSS.t272 17.4005
R3731 VSS.n439 VSS.t231 17.4005
R3732 VSS.n439 VSS.t226 17.4005
R3733 VSS.n442 VSS.t221 17.4005
R3734 VSS.n442 VSS.t277 17.4005
R3735 VSS.n443 VSS.t296 17.4005
R3736 VSS.n443 VSS.t233 17.4005
R3737 VSS.n446 VSS.t241 17.4005
R3738 VSS.n446 VSS.t239 17.4005
R3739 VSS.n447 VSS.t291 17.4005
R3740 VSS.n447 VSS.t289 17.4005
R3741 VSS.n450 VSS.t290 17.4005
R3742 VSS.n450 VSS.t245 17.4005
R3743 VSS.n451 VSS.t264 17.4005
R3744 VSS.n451 VSS.t293 17.4005
R3745 VSS.n869 VSS.t252 17.4005
R3746 VSS.n869 VSS.t230 17.4005
R3747 VSS.n870 VSS.t261 17.4005
R3748 VSS.n870 VSS.t247 17.4005
R3749 VSS.n872 VSS.t284 17.4005
R3750 VSS.n872 VSS.t286 17.4005
R3751 VSS.n873 VSS.t303 17.4005
R3752 VSS.n873 VSS.t283 17.4005
R3753 VSS.n875 VSS.t268 17.4005
R3754 VSS.n875 VSS.t243 17.4005
R3755 VSS.n877 VSS.t253 17.4005
R3756 VSS.n877 VSS.t228 17.4005
R3757 VSS.n878 VSS.t263 17.4005
R3758 VSS.n878 VSS.t250 17.4005
R3759 VSS.n880 VSS.t299 17.4005
R3760 VSS.n880 VSS.t298 17.4005
R3761 VSS.n882 VSS.t285 17.4005
R3762 VSS.n882 VSS.t287 17.4005
R3763 VSS.n883 VSS.t304 17.4005
R3764 VSS.n883 VSS.t281 17.4005
R3765 VSS.n885 VSS.t269 17.4005
R3766 VSS.n885 VSS.t244 17.4005
R3767 VSS.n887 VSS.t280 17.4005
R3768 VSS.n887 VSS.t257 17.4005
R3769 VSS.n888 VSS.t294 17.4005
R3770 VSS.n888 VSS.t279 17.4005
R3771 VSS.n890 VSS.t236 17.4005
R3772 VSS.n890 VSS.t232 17.4005
R3773 VSS.n892 VSS.t309 17.4005
R3774 VSS.n892 VSS.t310 17.4005
R3775 VSS.n893 VSS.t237 17.4005
R3776 VSS.n893 VSS.t308 17.4005
R3777 VSS.n895 VSS.t305 17.4005
R3778 VSS.n895 VSS.t271 17.4005
R3779 VSS.n897 VSS.t307 17.4005
R3780 VSS.n897 VSS.t288 17.4005
R3781 VSS.n898 VSS.t224 17.4005
R3782 VSS.n898 VSS.t306 17.4005
R3783 VSS.n900 VSS.t260 17.4005
R3784 VSS.n900 VSS.t258 17.4005
R3785 VSS.n902 VSS.t259 17.4005
R3786 VSS.n902 VSS.t238 17.4005
R3787 VSS.n903 VSS.t223 17.4005
R3788 VSS.n903 VSS.t300 17.4005
R3789 VSS.n906 VSS.t49 17.4005
R3790 VSS.n906 VSS.t103 17.4005
R3791 VSS.n923 VSS.t163 17.4005
R3792 VSS.n923 VSS.t157 17.4005
R3793 VSS.n916 VSS.t208 17.4005
R3794 VSS.n916 VSS.t90 17.4005
R3795 VSS.n913 VSS.t85 17.4005
R3796 VSS.n913 VSS.t72 17.4005
R3797 VSS.n3 VSS.t311 17.4005
R3798 VSS.n3 VSS.t251 17.4005
R3799 VSS.n4 VSS.t240 17.4005
R3800 VSS.n4 VSS.t267 17.4005
R3801 VSS.n6 VSS.t262 17.4005
R3802 VSS.n6 VSS.t295 17.4005
R3803 VSS.n49 VSS.t292 17.4005
R3804 VSS.n49 VSS.t210 17.4005
R3805 VSS.n45 VSS.t265 17.4005
R3806 VSS.n45 VSS.t173 17.4005
R3807 VSS.n38 VSS.t255 17.4005
R3808 VSS.n38 VSS.t143 17.4005
R3809 VSS.n33 VSS.t301 17.4005
R3810 VSS.n33 VSS.t31 17.4005
R3811 VSS.n27 VSS.t43 17.4005
R3812 VSS.n27 VSS.t254 17.4005
R3813 VSS.n94 VSS.t100 17.4005
R3814 VSS.n94 VSS.t270 17.4005
R3815 VSS.n19 VSS.t192 17.4005
R3816 VSS.n19 VSS.t227 17.4005
R3817 VSS.n104 VSS.t178 17.4005
R3818 VSS.n104 VSS.t220 17.4005
R3819 VSS.n112 VSS.t23 17.4005
R3820 VSS.n112 VSS.t242 17.4005
R3821 VSS.n115 VSS.t87 17.4005
R3822 VSS.n115 VSS.t248 17.4005
R3823 VSS.n84 VSS.t249 17.4005
R3824 VSS.n84 VSS.t282 17.4005
R3825 VSS.n82 VSS.t266 17.4005
R3826 VSS.n82 VSS.t302 17.4005
R3827 VSS.n81 VSS.t225 17.4005
R3828 VSS.n81 VSS.t256 17.4005
R3829 VSS.n78 VSS.t276 17.4005
R3830 VSS.n78 VSS.t184 17.4005
R3831 VSS.n43 VSS.t246 17.4005
R3832 VSS.n43 VSS.t134 17.4005
R3833 VSS.n1092 VSS.t198 17.4005
R3834 VSS.n1092 VSS.t46 17.4005
R3835 VSS.t46 VSS.n1091 17.4005
R3836 VSS.n1091 VSS.t36 17.4005
R3837 VSS.t182 VSS.n1024 17.4005
R3838 VSS.n1024 VSS.t176 17.4005
R3839 VSS.t150 VSS.n1025 17.4005
R3840 VSS.n1025 VSS.t182 17.4005
R3841 VSS.n1001 VSS.t204 17.4005
R3842 VSS.n1001 VSS.t167 17.4005
R3843 VSS.t167 VSS.n1000 17.4005
R3844 VSS.n1000 VSS.t169 17.4005
R3845 VSS.t130 VSS.n998 17.4005
R3846 VSS.n998 VSS.t69 17.4005
R3847 VSS.n993 VSS.t75 17.4005
R3848 VSS.n993 VSS.t78 17.4005
R3849 VSS.t169 VSS.n999 17.4005
R3850 VSS.n999 VSS.t130 17.4005
R3851 VSS.t78 VSS.n992 17.4005
R3852 VSS.n992 VSS.t159 17.4005
R3853 VSS.n1084 VSS.t112 17.4005
R3854 VSS.n1084 VSS.t118 17.4005
R3855 VSS.t36 VSS.n1090 17.4005
R3856 VSS.n1090 VSS.t96 17.4005
R3857 VSS.t96 VSS.n1089 17.4005
R3858 VSS.n1089 VSS.t25 17.4005
R3859 VSS.t118 VSS.n1083 17.4005
R3860 VSS.n1083 VSS.t189 17.4005
R3861 VSS.t82 VSS.n1006 17.4005
R3862 VSS.n1006 VSS.t120 17.4005
R3863 VSS.t120 VSS.n1005 17.4005
R3864 VSS.n1005 VSS.t116 17.4005
R3865 VSS.n501 VSS.n500 17.3498
R3866 VSS.n2385 VSS.n2384 17.3181
R3867 VSS.n1100 VSS.n1099 17.2121
R3868 VSS.n1224 VSS.t45 15.6539
R3869 VSS.n2358 VSS.t214 15.4735
R3870 VSS.n159 VSS.t219 15.4735
R3871 VSS.t13 VSS.n228 14.9582
R3872 VSS.n1285 VSS.t9 14.9582
R3873 VSS.n2158 VSS.t11 14.2625
R3874 VSS.n665 VSS.t48 14.2625
R3875 VSS.n1340 VSS.t8 14.2625
R3876 VSS.n1360 VSS.t77 14.2625
R3877 VSS.n1719 VSS.n1718 13.964
R3878 VSS.n2382 VSS.n125 13.964
R3879 VSS.n265 VSS.t156 13.5668
R3880 VSS.t212 VSS.n766 13.5668
R3881 VSS.n2387 VSS.n9 13.1961
R3882 VSS.n239 VSS.t7 12.8711
R3883 VSS.n656 VSS.n313 12.8711
R3884 VSS.n1243 VSS.t16 12.8711
R3885 VSS.n1718 VSS.n125 11.6996
R3886 VSS.n810 VSS.t16 10.784
R3887 VSS.n2097 VSS.n667 10.5417
R3888 VSS.n953 VSS.n952 10.4392
R3889 VSS.n152 VSS.t214 10.1901
R3890 VSS.n2350 VSS.t219 10.1901
R3891 VSS.t7 VSS.n235 10.0883
R3892 VSS.n1297 VSS.t212 10.0883
R3893 VSS.n645 VSS.t14 9.39255
R3894 VSS.n655 VSS.t213 9.39255
R3895 VSS.n2122 VSS.t48 9.39255
R3896 VSS.n1347 VSS.t8 9.39255
R3897 VSS.n1353 VSS.t77 9.39255
R3898 VSS.n952 VSS.n667 9.3005
R3899 VSS.n2386 VSS.n2385 9.3005
R3900 VSS.n2131 VSS.n313 9.04469
R3901 VSS.n2203 VSS.t13 8.69684
R3902 VSS.n2187 VSS.t162 8.69684
R3903 VSS.t9 VSS.n774 8.69684
R3904 VSS.n499 VSS.n498 8.69572
R3905 VSS.n1783 VSS.n1618 8.35212
R3906 VSS.n498 VSS.n497 8.00322
R3907 VSS.t18 VSS.t162 8.00113
R3908 VSS.t156 VSS.t0 8.00113
R3909 VSS.t14 VSS.t312 8.00113
R3910 VSS.t213 VSS.t51 8.00113
R3911 VSS.n1231 VSS.t45 8.00113
R3912 VSS.n1099 VSS.n1098 7.97904
R3913 VSS.n2392 VSS.n2391 7.91206
R3914 VSS.n637 VSS.t11 7.65328
R3915 VSS.n1782 VSS.n1781 6.41614
R3916 VSS.n1101 VSS.n1100 6.4005
R3917 VSS.n938 VSS.n937 6.34833
R3918 VSS.n802 VSS.t15 5.91401
R3919 VSS.n87 VSS.n86 5.74088
R3920 VSS.n86 VSS.n80 5.74088
R3921 VSS.t22 VSS.n126 5.66136
R3922 VSS.n1087 VSS.n1086 5.46789
R3923 VSS.n1047 VSS.n1046 5.46789
R3924 VSS.n615 VSS.t18 5.2183
R3925 VSS.n1309 VSS.t19 5.2183
R3926 VSS.n1780 VSS.n1717 4.90658
R3927 VSS.n145 VSS.t215 4.90658
R3928 VSS.n2342 VSS.t30 4.90658
R3929 VSS.n86 VSS.n85 4.5872
R3930 VSS.n2145 VSS.t312 4.5226
R3931 VSS.t51 VSS.n307 4.5226
R3932 VSS.n2114 VSS.t102 4.5226
R3933 VSS.n1334 VSS.t12 4.5226
R3934 VSS.n1367 VSS.t38 4.5226
R3935 VSS.n1210 VSS.n1208 4.17474
R3936 VSS.n1209 VSS.n821 4.17474
R3937 VSS.n822 VSS.n817 4.17474
R3938 VSS.n1225 VSS.n1223 4.17474
R3939 VSS.n2211 VSS.t10 3.82689
R3940 VSS.n2123 VSS.n2122 3.82689
R3941 VSS.t6 VSS.n782 3.82689
R3942 VSS.n2166 VSS.t313 3.47904
R3943 VSS.t56 VSS.n1216 3.13118
R3944 VSS.n961 VSS.n0 2.83186
R3945 VSS.t1 VSS.n274 2.78333
R3946 VSS VSS.n2392 2.40512
R3947 VSS.n1785 VSS.n1784 2.17107
R3948 VSS.n1778 VSS.n1777 2.17107
R3949 VSS.n1777 VSS.n1776 2.17107
R3950 VSS.n2003 VSS.t4 1.75629
R3951 VSS.n2193 VSS.n242 1.73977
R3952 VSS.n615 VSS.n614 1.73977
R3953 VSS.n2187 VSS.n2186 1.73977
R3954 VSS.n619 VSS.n249 1.73977
R3955 VSS.n2180 VSS.n257 1.73977
R3956 VSS.n2179 VSS.n259 1.73977
R3957 VSS.n266 VSS.n265 1.73977
R3958 VSS.n2173 VSS.n2172 1.73977
R3959 VSS.n628 VSS.n268 1.73977
R3960 VSS.n2166 VSS.n274 1.73977
R3961 VSS.n2165 VSS.n276 1.73977
R3962 VSS.n283 VSS.n282 1.73977
R3963 VSS.n2159 VSS.n2158 1.73977
R3964 VSS.n2152 VSS.n290 1.73977
R3965 VSS.n2151 VSS.n292 1.73977
R3966 VSS.n645 VSS.n644 1.73977
R3967 VSS.n2145 VSS.n2144 1.73977
R3968 VSS.n649 VSS.n299 1.73977
R3969 VSS.n2138 VSS.n305 1.73977
R3970 VSS.n2137 VSS.n307 1.73977
R3971 VSS.n656 VSS.n655 1.73977
R3972 VSS.n2131 VSS.n2130 1.73977
R3973 VSS.n1778 VSS.n9 1.62843
R3974 VSS.n960 VSS.n871 1.56325
R3975 VSS.n2389 VSS.n7 1.5223
R3976 VSS.n2389 VSS.n2388 1.40267
R3977 VSS.n2390 VSS.n2389 1.40267
R3978 VSS.n638 VSS.t217 1.39191
R3979 VSS.n959 VSS.n876 1.22642
R3980 VSS.n957 VSS.n886 1.22642
R3981 VSS.n955 VSS.n896 1.22642
R3982 VSS.n953 VSS.n904 1.22642
R3983 VSS.n1097 VSS.n963 1.18528
R3984 VSS.n976 VSS.n972 1.18528
R3985 VSS.n2392 VSS.n0 1.16343
R3986 VSS.n7 VSS.n5 1.1365
R3987 VSS.n1056 VSS.n1055 1.13093
R3988 VSS.n1045 VSS.n1044 1.13093
R3989 VSS.n589 VSS.n501 1.12991
R3990 VSS.n85 VSS.n83 1.10524
R3991 VSS.n2219 VSS.t27 1.04406
R3992 VSS.n1217 VSS.t56 1.04406
R3993 VSS.n794 VSS.t17 1.04406
R3994 VSS.n2388 VSS.n8 1.03854
R3995 VSS.n2390 VSS.n2 1.03854
R3996 VSS.n1088 VSS.n1087 0.911718
R3997 VSS.n1086 VSS.n1085 0.911718
R3998 VSS.n969 VSS.n968 0.911718
R3999 VSS.n2391 VSS.n1 0.891397
R4000 VSS.n958 VSS.n881 0.889583
R4001 VSS.n956 VSS.n891 0.889583
R4002 VSS.n954 VSS.n901 0.889583
R4003 VSS.n437 VSS.n436 0.886319
R4004 VSS.n445 VSS.n444 0.886319
R4005 VSS.n453 VSS.n452 0.886319
R4006 VSS.n2387 VSS.n2386 0.82387
R4007 VSS.n437 VSS.n433 0.775347
R4008 VSS.n2391 VSS.n2390 0.739223
R4009 VSS.n106 VSS.n105 0.709873
R4010 VSS.n88 VSS.n25 0.709873
R4011 VSS.n31 VSS.n29 0.709873
R4012 VSS.n44 VSS.n41 0.709873
R4013 VSS.n925 VSS.n922 0.709871
R4014 VSS.n99 VSS.n20 0.709871
R4015 VSS.n68 VSS.n39 0.709871
R4016 VSS.n1062 VSS.n986 0.709871
R4017 VSS.n2388 VSS.n2387 0.701587
R4018 VSS.n2195 VSS.n239 0.696207
R4019 VSS.n876 VSS.n874 0.674167
R4020 VSS.n881 VSS.n879 0.674167
R4021 VSS.n886 VSS.n884 0.674167
R4022 VSS.n891 VSS.n889 0.674167
R4023 VSS.n896 VSS.n894 0.674167
R4024 VSS.n901 VSS.n899 0.674167
R4025 VSS.n969 VSS.n963 0.630935
R4026 VSS.n1047 VSS.n991 0.630935
R4027 VSS.n1054 VSS.n991 0.630935
R4028 VSS.n970 VSS.n969 0.630935
R4029 VSS.n1087 VSS.n970 0.630935
R4030 VSS.n1086 VSS.n972 0.630935
R4031 VSS.n1055 VSS.n1054 0.630935
R4032 VSS.n1046 VSS.n1045 0.630935
R4033 VSS.n88 VSS.n87 0.591912
R4034 VSS.n80 VSS.n29 0.591912
R4035 VSS.n996 VSS.n995 0.570371
R4036 VSS.n1023 VSS.n1022 0.570371
R4037 VSS.n441 VSS.n440 0.549486
R4038 VSS.n449 VSS.n448 0.549486
R4039 VSS.n1784 VSS.n9 0.543143
R4040 VSS.n1081 VSS.n972 0.484196
R4041 VSS.n964 VSS.n963 0.484196
R4042 VSS.n1099 VSS.n961 0.43055
R4043 VSS.n1054 VSS.n1053 0.428385
R4044 VSS.n1048 VSS.n1047 0.428385
R4045 VSS.n1046 VSS.n1002 0.428385
R4046 VSS.n1050 VSS.n991 0.421696
R4047 VSS.n1055 VSS.n990 0.421696
R4048 VSS.n1045 VSS.n1004 0.421696
R4049 VSS.t216 VSS.n135 0.377891
R4050 VSS.n927 VSS.n921 0.367414
R4051 VSS.n929 VSS.n920 0.367414
R4052 VSS.n931 VSS.n919 0.367414
R4053 VSS.n935 VSS.n915 0.367414
R4054 VSS.n484 VSS.n482 0.359263
R4055 VSS.n486 VSS.n481 0.359263
R4056 VSS.n488 VSS.n480 0.359263
R4057 VSS.n490 VSS.n479 0.359263
R4058 VSS.n492 VSS.n478 0.359263
R4059 VSS.n494 VSS.n477 0.359263
R4060 VSS.n496 VSS.n476 0.359263
R4061 VSS.n462 VSS.n460 0.359263
R4062 VSS.n464 VSS.n459 0.359263
R4063 VSS.n466 VSS.n458 0.359263
R4064 VSS.n468 VSS.n457 0.359263
R4065 VSS.n470 VSS.n456 0.359263
R4066 VSS.n472 VSS.n455 0.359263
R4067 VSS.n474 VSS.n454 0.359263
R4068 VSS.n926 VSS.n922 0.359263
R4069 VSS.n928 VSS.n921 0.359263
R4070 VSS.n930 VSS.n920 0.359263
R4071 VSS.n932 VSS.n919 0.359263
R4072 VSS.n934 VSS.n918 0.359263
R4073 VSS.n937 VSS.n915 0.359263
R4074 VSS.n938 VSS.n912 0.359263
R4075 VSS.n941 VSS.n911 0.359263
R4076 VSS.n943 VSS.n910 0.359263
R4077 VSS.n945 VSS.n909 0.359263
R4078 VSS.n947 VSS.n908 0.359263
R4079 VSS.n949 VSS.n905 0.359263
R4080 VSS.n11 VSS.n10 0.359263
R4081 VSS.n117 VSS.n116 0.359263
R4082 VSS.n111 VSS.n109 0.359263
R4083 VSS.n113 VSS.n13 0.359263
R4084 VSS.n103 VSS.n15 0.359263
R4085 VSS.n101 VSS.n17 0.359263
R4086 VSS.n21 VSS.n18 0.359263
R4087 VSS.n97 VSS.n20 0.359263
R4088 VSS.n93 VSS.n91 0.359263
R4089 VSS.n95 VSS.n23 0.359263
R4090 VSS.n74 VSS.n32 0.359263
R4091 VSS.n34 VSS.n30 0.359263
R4092 VSS.n70 VSS.n36 0.359263
R4093 VSS.n39 VSS.n37 0.359263
R4094 VSS.n66 VSS.n40 0.359263
R4095 VSS.n64 VSS.n63 0.359263
R4096 VSS.n59 VSS.n46 0.359263
R4097 VSS.n48 VSS.n42 0.359263
R4098 VSS.n51 VSS.n50 0.359263
R4099 VSS.n55 VSS.n54 0.359263
R4100 VSS.n1078 VSS.n977 0.359263
R4101 VSS.n1076 VSS.n978 0.359263
R4102 VSS.n1074 VSS.n979 0.359263
R4103 VSS.n1072 VSS.n980 0.359263
R4104 VSS.n1070 VSS.n981 0.359263
R4105 VSS.n1068 VSS.n982 0.359263
R4106 VSS.n1066 VSS.n983 0.359263
R4107 VSS.n1064 VSS.n984 0.359263
R4108 VSS.n1060 VSS.n985 0.359263
R4109 VSS.n1056 VSS.n988 0.359263
R4110 VSS.n1044 VSS.n1007 0.359263
R4111 VSS.n1041 VSS.n1008 0.359263
R4112 VSS.n1039 VSS.n1009 0.359263
R4113 VSS.n1037 VSS.n1010 0.359263
R4114 VSS.n1035 VSS.n1011 0.359263
R4115 VSS.n1033 VSS.n1012 0.359263
R4116 VSS.n1031 VSS.n1013 0.359263
R4117 VSS.n1029 VSS.n1014 0.359263
R4118 VSS.n1027 VSS.n1026 0.359263
R4119 VSS.n485 VSS.n482 0.359261
R4120 VSS.n487 VSS.n481 0.359261
R4121 VSS.n489 VSS.n480 0.359261
R4122 VSS.n491 VSS.n479 0.359261
R4123 VSS.n493 VSS.n478 0.359261
R4124 VSS.n495 VSS.n477 0.359261
R4125 VSS.n497 VSS.n476 0.359261
R4126 VSS.n463 VSS.n460 0.359261
R4127 VSS.n465 VSS.n459 0.359261
R4128 VSS.n467 VSS.n458 0.359261
R4129 VSS.n469 VSS.n457 0.359261
R4130 VSS.n471 VSS.n456 0.359261
R4131 VSS.n473 VSS.n455 0.359261
R4132 VSS.n475 VSS.n454 0.359261
R4133 VSS.n933 VSS.n918 0.359261
R4134 VSS.n940 VSS.n912 0.359261
R4135 VSS.n942 VSS.n911 0.359261
R4136 VSS.n944 VSS.n910 0.359261
R4137 VSS.n946 VSS.n909 0.359261
R4138 VSS.n948 VSS.n908 0.359261
R4139 VSS.n951 VSS.n905 0.359261
R4140 VSS.n120 VSS.n10 0.359261
R4141 VSS.n116 VSS.n8 0.359261
R4142 VSS.n111 VSS.n110 0.359261
R4143 VSS.n114 VSS.n113 0.359261
R4144 VSS.n108 VSS.n15 0.359261
R4145 VSS.n105 VSS.n16 0.359261
R4146 VSS.n102 VSS.n17 0.359261
R4147 VSS.n100 VSS.n18 0.359261
R4148 VSS.n93 VSS.n92 0.359261
R4149 VSS.n96 VSS.n95 0.359261
R4150 VSS.n90 VSS.n25 0.359261
R4151 VSS.n75 VSS.n31 0.359261
R4152 VSS.n71 VSS.n32 0.359261
R4153 VSS.n35 VSS.n34 0.359261
R4154 VSS.n67 VSS.n36 0.359261
R4155 VSS.n65 VSS.n40 0.359261
R4156 VSS.n60 VSS.n44 0.359261
R4157 VSS.n63 VSS.n62 0.359261
R4158 VSS.n47 VSS.n46 0.359261
R4159 VSS.n56 VSS.n48 0.359261
R4160 VSS.n50 VSS.n2 0.359261
R4161 VSS.n54 VSS.n1 0.359261
R4162 VSS.n977 VSS.n976 0.359261
R4163 VSS.n1082 VSS.n1081 0.359261
R4164 VSS.n1077 VSS.n978 0.359261
R4165 VSS.n1075 VSS.n979 0.359261
R4166 VSS.n1073 VSS.n980 0.359261
R4167 VSS.n1071 VSS.n981 0.359261
R4168 VSS.n1069 VSS.n982 0.359261
R4169 VSS.n1067 VSS.n983 0.359261
R4170 VSS.n1065 VSS.n984 0.359261
R4171 VSS.n1063 VSS.n985 0.359261
R4172 VSS.n1059 VSS.n988 0.359261
R4173 VSS.n997 VSS.n989 0.359261
R4174 VSS.n1042 VSS.n1007 0.359261
R4175 VSS.n1040 VSS.n1008 0.359261
R4176 VSS.n1038 VSS.n1009 0.359261
R4177 VSS.n1036 VSS.n1010 0.359261
R4178 VSS.n1034 VSS.n1011 0.359261
R4179 VSS.n1032 VSS.n1012 0.359261
R4180 VSS.n1030 VSS.n1013 0.359261
R4181 VSS.n1028 VSS.n1014 0.359261
R4182 VSS.n1026 VSS.n1017 0.359261
R4183 VSS.n1018 VSS.n966 0.359261
R4184 VSS.n1093 VSS.n964 0.359261
R4185 VSS.n965 VSS.n962 0.357865
R4186 VSS.n1082 VSS.n975 0.351111
R4187 VSS.n987 VSS.n986 0.351111
R4188 VSS.n997 VSS.n990 0.351111
R4189 VSS.n1019 VSS.n1018 0.351111
R4190 VSS.n1094 VSS.n1093 0.351111
R4191 VSS.n925 VSS.n924 0.35111
R4192 VSS.n937 VSS.n936 0.35111
R4193 VSS.n936 VSS.n917 0.35111
R4194 VSS.n939 VSS.n914 0.35111
R4195 VSS.n939 VSS.n938 0.35111
R4196 VSS.n950 VSS.n907 0.35111
R4197 VSS.n951 VSS.n950 0.35111
R4198 VSS.n120 VSS.n119 0.35111
R4199 VSS.n119 VSS.n8 0.35111
R4200 VSS.n118 VSS.n11 0.35111
R4201 VSS.n118 VSS.n117 0.35111
R4202 VSS.n110 VSS.n12 0.35111
R4203 VSS.n114 VSS.n12 0.35111
R4204 VSS.n109 VSS.n14 0.35111
R4205 VSS.n14 VSS.n13 0.35111
R4206 VSS.n108 VSS.n107 0.35111
R4207 VSS.n107 VSS.n16 0.35111
R4208 VSS.n106 VSS.n103 0.35111
R4209 VSS.n100 VSS.n99 0.35111
R4210 VSS.n98 VSS.n21 0.35111
R4211 VSS.n98 VSS.n97 0.35111
R4212 VSS.n92 VSS.n22 0.35111
R4213 VSS.n96 VSS.n22 0.35111
R4214 VSS.n91 VSS.n24 0.35111
R4215 VSS.n24 VSS.n23 0.35111
R4216 VSS.n90 VSS.n89 0.35111
R4217 VSS.n89 VSS.n26 0.35111
R4218 VSS.n77 VSS.n76 0.35111
R4219 VSS.n76 VSS.n75 0.35111
R4220 VSS.n73 VSS.n30 0.35111
R4221 VSS.n74 VSS.n73 0.35111
R4222 VSS.n72 VSS.n35 0.35111
R4223 VSS.n72 VSS.n71 0.35111
R4224 VSS.n69 VSS.n37 0.35111
R4225 VSS.n70 VSS.n69 0.35111
R4226 VSS.n68 VSS.n67 0.35111
R4227 VSS.n64 VSS.n41 0.35111
R4228 VSS.n61 VSS.n60 0.35111
R4229 VSS.n62 VSS.n61 0.35111
R4230 VSS.n59 VSS.n58 0.35111
R4231 VSS.n58 VSS.n42 0.35111
R4232 VSS.n57 VSS.n47 0.35111
R4233 VSS.n57 VSS.n56 0.35111
R4234 VSS.n53 VSS.n51 0.35111
R4235 VSS.n55 VSS.n53 0.35111
R4236 VSS.n52 VSS.n2 0.35111
R4237 VSS.n52 VSS.n1 0.35111
R4238 VSS.n1095 VSS.n965 0.35111
R4239 VSS.n1081 VSS.n1080 0.35111
R4240 VSS.n1080 VSS.n976 0.35111
R4241 VSS.n1079 VSS.n1078 0.35111
R4242 VSS.n1063 VSS.n1062 0.35111
R4243 VSS.n1061 VSS.n1060 0.35111
R4244 VSS.n1058 VSS.n989 0.35111
R4245 VSS.n1059 VSS.n1058 0.35111
R4246 VSS.n1057 VSS.n1056 0.35111
R4247 VSS.n1044 VSS.n1043 0.35111
R4248 VSS.n1027 VSS.n1015 0.35111
R4249 VSS.n1017 VSS.n1016 0.35111
R4250 VSS.n1016 VSS.n966 0.35111
R4251 VSS.n1097 VSS.n1096 0.35111
R4252 VSS.n1096 VSS.n964 0.35111
R4253 VSS.t0 VSS.n259 0.348354
R4254 VSS.t217 VSS.n637 0.348354
R4255 VSS.n1321 VSS.t20 0.348354
R4256 VSS.n484 VSS.n483 0.3483
R4257 VSS.n462 VSS.n461 0.3483
R4258 VSS.n1095 VSS.n1094 0.343898
R4259 VSS.n1079 VSS.n975 0.343898
R4260 VSS.n1061 VSS.n987 0.343898
R4261 VSS.n1057 VSS.n990 0.343898
R4262 VSS.n1043 VSS.n1004 0.343898
R4263 VSS.n1019 VSS.n1015 0.343898
R4264 VSS.n28 VSS.n26 0.328001
R4265 VSS.n79 VSS.n77 0.328001
R4266 VSS.n1053 VSS.n996 0.310758
R4267 VSS.n1088 VSS.n971 0.310758
R4268 VSS.n1085 VSS.n973 0.310758
R4269 VSS.n1023 VSS.n1021 0.310758
R4270 VSS.n1022 VSS.n968 0.310758
R4271 VSS.n974 VSS.n973 0.310756
R4272 VSS.n975 VSS.n974 0.310756
R4273 VSS.n995 VSS.n994 0.310756
R4274 VSS.n994 VSS.n987 0.310756
R4275 VSS.n1049 VSS.n1048 0.310756
R4276 VSS.n1050 VSS.n1049 0.310756
R4277 VSS.n1051 VSS.n1050 0.310756
R4278 VSS.n1053 VSS.n1051 0.310756
R4279 VSS.n1053 VSS.n1052 0.310756
R4280 VSS.n1052 VSS.n990 0.310756
R4281 VSS.n1004 VSS.n1003 0.310756
R4282 VSS.n1003 VSS.n1002 0.310756
R4283 VSS.n1020 VSS.n1019 0.310756
R4284 VSS.n1021 VSS.n1020 0.310756
R4285 VSS.n1094 VSS.n967 0.310756
R4286 VSS.n1022 VSS.n967 0.310756
R4287 VSS.n952 VSS.n951 0.310283
R4288 VSS.n498 VSS.n475 0.291261
R4289 VSS.n441 VSS.n437 0.226361
R4290 VSS.n445 VSS.n441 0.226361
R4291 VSS.n449 VSS.n445 0.226361
R4292 VSS.n453 VSS.n449 0.226361
R4293 VSS.n500 VSS.n453 0.226361
R4294 VSS.n960 VSS.n959 0.226361
R4295 VSS.n959 VSS.n958 0.226361
R4296 VSS.n958 VSS.n957 0.226361
R4297 VSS.n957 VSS.n956 0.226361
R4298 VSS.n956 VSS.n955 0.226361
R4299 VSS.n955 VSS.n954 0.226361
R4300 VSS.n954 VSS.n953 0.226361
R4301 VSS.n961 VSS.n960 0.222444
R4302 VSS.n2386 VSS.n120 0.215174
R4303 VSS.n947 VSS.n946 0.179848
R4304 VSS.n949 VSS.n948 0.179848
R4305 VSS.n1098 VSS.n1097 0.174309
R4306 VSS.n927 VSS.n926 0.171696
R4307 VSS.n929 VSS.n928 0.171696
R4308 VSS.n486 VSS.n485 0.168978
R4309 VSS.n488 VSS.n487 0.168978
R4310 VSS.n490 VSS.n489 0.168978
R4311 VSS.n492 VSS.n491 0.168978
R4312 VSS.n494 VSS.n493 0.168978
R4313 VSS.n496 VSS.n495 0.168978
R4314 VSS.n464 VSS.n463 0.168978
R4315 VSS.n466 VSS.n465 0.168978
R4316 VSS.n468 VSS.n467 0.168978
R4317 VSS.n470 VSS.n469 0.168978
R4318 VSS.n472 VSS.n471 0.168978
R4319 VSS.n474 VSS.n473 0.168978
R4320 VSS.n933 VSS.n932 0.168978
R4321 VSS.n941 VSS.n940 0.168978
R4322 VSS.n943 VSS.n942 0.168978
R4323 VSS.n945 VSS.n944 0.168978
R4324 VSS.n117 VSS.n114 0.168978
R4325 VSS.n110 VSS.n11 0.168978
R4326 VSS.n16 VSS.n13 0.168978
R4327 VSS.n109 VSS.n108 0.168978
R4328 VSS.n103 VSS.n102 0.168978
R4329 VSS.n101 VSS.n100 0.168978
R4330 VSS.n97 VSS.n96 0.168978
R4331 VSS.n92 VSS.n21 0.168978
R4332 VSS.n26 VSS.n23 0.168978
R4333 VSS.n91 VSS.n90 0.168978
R4334 VSS.n77 VSS.n30 0.168978
R4335 VSS.n75 VSS.n74 0.168978
R4336 VSS.n37 VSS.n35 0.168978
R4337 VSS.n71 VSS.n70 0.168978
R4338 VSS.n67 VSS.n66 0.168978
R4339 VSS.n65 VSS.n64 0.168978
R4340 VSS.n62 VSS.n42 0.168978
R4341 VSS.n60 VSS.n59 0.168978
R4342 VSS.n56 VSS.n55 0.168978
R4343 VSS.n51 VSS.n47 0.168978
R4344 VSS.n1078 VSS.n1077 0.168978
R4345 VSS.n1076 VSS.n1075 0.168978
R4346 VSS.n1074 VSS.n1073 0.168978
R4347 VSS.n1072 VSS.n1071 0.168978
R4348 VSS.n1070 VSS.n1069 0.168978
R4349 VSS.n1068 VSS.n1067 0.168978
R4350 VSS.n1066 VSS.n1065 0.168978
R4351 VSS.n1064 VSS.n1063 0.168978
R4352 VSS.n1060 VSS.n1059 0.168978
R4353 VSS.n1042 VSS.n1041 0.168978
R4354 VSS.n1040 VSS.n1039 0.168978
R4355 VSS.n1038 VSS.n1037 0.168978
R4356 VSS.n1036 VSS.n1035 0.168978
R4357 VSS.n1034 VSS.n1033 0.168978
R4358 VSS.n1032 VSS.n1031 0.168978
R4359 VSS.n1030 VSS.n1029 0.168978
R4360 VSS.n1028 VSS.n1027 0.168978
R4361 VSS.n1017 VSS.n965 0.168978
R4362 VSS.n1098 VSS.n962 0.164301
R4363 VSS.n931 VSS.n930 0.160826
R4364 VSS.n935 VSS.n934 0.160826
R4365 VSS.n1094 VSS.n966 0.160826
R4366 VSS.n989 VSS.n987 0.160826
R4367 VSS.n500 VSS.n499 0.136278
R4368 VSS.n499 VSS.n0 0.109514
R4369 VSS.n87 VSS.n28 0.0871999
R4370 VSS.n80 VSS.n79 0.0871999
R4371 a_8862_4192.n21 a_8862_4192.n19 70.8255
R4372 a_8862_4192.n2 a_8862_4192.n0 70.8255
R4373 a_8862_4192.n14 a_8862_4192.n13 69.6895
R4374 a_8862_4192.n16 a_8862_4192.n15 69.6895
R4375 a_8862_4192.n18 a_8862_4192.n17 69.6895
R4376 a_8862_4192.n23 a_8862_4192.n22 69.6895
R4377 a_8862_4192.n21 a_8862_4192.n20 69.6895
R4378 a_8862_4192.n12 a_8862_4192.n11 69.6895
R4379 a_8862_4192.n10 a_8862_4192.n9 69.6895
R4380 a_8862_4192.n8 a_8862_4192.n7 69.6895
R4381 a_8862_4192.n6 a_8862_4192.n5 69.6895
R4382 a_8862_4192.n4 a_8862_4192.n3 69.6895
R4383 a_8862_4192.n2 a_8862_4192.n1 69.6895
R4384 a_8862_4192.n25 a_8862_4192.n24 69.6895
R4385 a_8862_4192.n13 a_8862_4192.t22 17.4005
R4386 a_8862_4192.n13 a_8862_4192.t21 17.4005
R4387 a_8862_4192.n15 a_8862_4192.t26 17.4005
R4388 a_8862_4192.n15 a_8862_4192.t25 17.4005
R4389 a_8862_4192.n17 a_8862_4192.t14 17.4005
R4390 a_8862_4192.n17 a_8862_4192.t13 17.4005
R4391 a_8862_4192.n22 a_8862_4192.t11 17.4005
R4392 a_8862_4192.n22 a_8862_4192.t9 17.4005
R4393 a_8862_4192.n20 a_8862_4192.t19 17.4005
R4394 a_8862_4192.n20 a_8862_4192.t17 17.4005
R4395 a_8862_4192.n19 a_8862_4192.t24 17.4005
R4396 a_8862_4192.n19 a_8862_4192.t23 17.4005
R4397 a_8862_4192.n11 a_8862_4192.t12 17.4005
R4398 a_8862_4192.n11 a_8862_4192.t10 17.4005
R4399 a_8862_4192.n9 a_8862_4192.t20 17.4005
R4400 a_8862_4192.n9 a_8862_4192.t18 17.4005
R4401 a_8862_4192.n7 a_8862_4192.t6 17.4005
R4402 a_8862_4192.n7 a_8862_4192.t5 17.4005
R4403 a_8862_4192.n5 a_8862_4192.t2 17.4005
R4404 a_8862_4192.n5 a_8862_4192.t1 17.4005
R4405 a_8862_4192.n3 a_8862_4192.t4 17.4005
R4406 a_8862_4192.n3 a_8862_4192.t27 17.4005
R4407 a_8862_4192.n1 a_8862_4192.t8 17.4005
R4408 a_8862_4192.n1 a_8862_4192.t7 17.4005
R4409 a_8862_4192.n0 a_8862_4192.t16 17.4005
R4410 a_8862_4192.n0 a_8862_4192.t15 17.4005
R4411 a_8862_4192.t0 a_8862_4192.n25 17.4005
R4412 a_8862_4192.n25 a_8862_4192.t3 17.4005
R4413 a_8862_4192.n14 a_8862_4192.n12 3.84846
R4414 a_8862_4192.n16 a_8862_4192.n14 1.1365
R4415 a_8862_4192.n12 a_8862_4192.n10 1.1365
R4416 a_8862_4192.n10 a_8862_4192.n8 1.1365
R4417 a_8862_4192.n8 a_8862_4192.n6 1.1365
R4418 a_8862_4192.n6 a_8862_4192.n4 1.1365
R4419 a_8862_4192.n4 a_8862_4192.n2 1.1365
R4420 a_8862_4192.n18 a_8862_4192.n16 1.1365
R4421 a_8862_4192.n24 a_8862_4192.n18 1.1365
R4422 a_8862_4192.n24 a_8862_4192.n23 1.1365
R4423 a_8862_4192.n23 a_8862_4192.n21 1.1365
R4424 VDD.n799 VDD.n557 758.823
R4425 VDD.n364 VDD.n98 758.823
R4426 VDD.n120 VDD.n96 758.823
R4427 VDD.n796 VDD.n572 702.354
R4428 VDD.n722 VDD.n657 660
R4429 VDD.n151 VDD.n125 660
R4430 VDD.n237 VDD.n127 660
R4431 VDD.n720 VDD.n659 603.529
R4432 VDD.n722 VDD.n655 240
R4433 VDD.n726 VDD.n655 240
R4434 VDD.n726 VDD.n649 240
R4435 VDD.n734 VDD.n649 240
R4436 VDD.n734 VDD.n647 240
R4437 VDD.n738 VDD.n647 240
R4438 VDD.n738 VDD.n641 240
R4439 VDD.n747 VDD.n641 240
R4440 VDD.n747 VDD.n639 240
R4441 VDD.n751 VDD.n639 240
R4442 VDD.n751 VDD.n634 240
R4443 VDD.n760 VDD.n634 240
R4444 VDD.n760 VDD.n632 240
R4445 VDD.n764 VDD.n632 240
R4446 VDD.n764 VDD.n627 240
R4447 VDD.n773 VDD.n627 240
R4448 VDD.n773 VDD.n625 240
R4449 VDD.n777 VDD.n625 240
R4450 VDD.n777 VDD.n620 240
R4451 VDD.n786 VDD.n620 240
R4452 VDD.n786 VDD.n618 240
R4453 VDD.n790 VDD.n618 240
R4454 VDD.n790 VDD.n557 240
R4455 VDD.n672 VDD.n657 240
R4456 VDD.n676 VDD.n674 240
R4457 VDD.n680 VDD.n669 240
R4458 VDD.n684 VDD.n682 240
R4459 VDD.n688 VDD.n667 240
R4460 VDD.n692 VDD.n690 240
R4461 VDD.n696 VDD.n665 240
R4462 VDD.n700 VDD.n698 240
R4463 VDD.n704 VDD.n663 240
R4464 VDD.n708 VDD.n706 240
R4465 VDD.n712 VDD.n661 240
R4466 VDD.n716 VDD.n714 240
R4467 VDD.n720 VDD.n653 240
R4468 VDD.n728 VDD.n653 240
R4469 VDD.n728 VDD.n651 240
R4470 VDD.n732 VDD.n651 240
R4471 VDD.n732 VDD.n645 240
R4472 VDD.n740 VDD.n645 240
R4473 VDD.n740 VDD.n643 240
R4474 VDD.n744 VDD.n643 240
R4475 VDD.n744 VDD.n638 240
R4476 VDD.n753 VDD.n638 240
R4477 VDD.n753 VDD.n636 240
R4478 VDD.n757 VDD.n636 240
R4479 VDD.n757 VDD.n631 240
R4480 VDD.n766 VDD.n631 240
R4481 VDD.n766 VDD.n629 240
R4482 VDD.n770 VDD.n629 240
R4483 VDD.n770 VDD.n624 240
R4484 VDD.n779 VDD.n624 240
R4485 VDD.n779 VDD.n622 240
R4486 VDD.n783 VDD.n622 240
R4487 VDD.n783 VDD.n617 240
R4488 VDD.n792 VDD.n617 240
R4489 VDD.n792 VDD.n572 240
R4490 VDD.n799 VDD.n558 240
R4491 VDD.n575 VDD.n574 240
R4492 VDD.n579 VDD.n578 240
R4493 VDD.n583 VDD.n582 240
R4494 VDD.n587 VDD.n586 240
R4495 VDD.n591 VDD.n590 240
R4496 VDD.n595 VDD.n594 240
R4497 VDD.n599 VDD.n598 240
R4498 VDD.n603 VDD.n602 240
R4499 VDD.n607 VDD.n606 240
R4500 VDD.n611 VDD.n610 240
R4501 VDD.n613 VDD.n571 240
R4502 VDD.n245 VDD.n125 240
R4503 VDD.n245 VDD.n123 240
R4504 VDD.n249 VDD.n123 240
R4505 VDD.n249 VDD.n63 240
R4506 VDD.n400 VDD.n63 240
R4507 VDD.n400 VDD.n64 240
R4508 VDD.n396 VDD.n64 240
R4509 VDD.n396 VDD.n70 240
R4510 VDD.n392 VDD.n70 240
R4511 VDD.n392 VDD.n72 240
R4512 VDD.n388 VDD.n72 240
R4513 VDD.n388 VDD.n77 240
R4514 VDD.n384 VDD.n77 240
R4515 VDD.n384 VDD.n79 240
R4516 VDD.n380 VDD.n79 240
R4517 VDD.n380 VDD.n84 240
R4518 VDD.n376 VDD.n84 240
R4519 VDD.n376 VDD.n86 240
R4520 VDD.n372 VDD.n86 240
R4521 VDD.n372 VDD.n91 240
R4522 VDD.n368 VDD.n91 240
R4523 VDD.n368 VDD.n93 240
R4524 VDD.n364 VDD.n93 240
R4525 VDD.n155 VDD.n154 240
R4526 VDD.n159 VDD.n158 240
R4527 VDD.n163 VDD.n162 240
R4528 VDD.n167 VDD.n166 240
R4529 VDD.n171 VDD.n170 240
R4530 VDD.n175 VDD.n174 240
R4531 VDD.n179 VDD.n178 240
R4532 VDD.n183 VDD.n182 240
R4533 VDD.n187 VDD.n186 240
R4534 VDD.n191 VDD.n190 240
R4535 VDD.n195 VDD.n194 240
R4536 VDD.n199 VDD.n198 240
R4537 VDD.n203 VDD.n202 240
R4538 VDD.n207 VDD.n206 240
R4539 VDD.n211 VDD.n210 240
R4540 VDD.n215 VDD.n214 240
R4541 VDD.n219 VDD.n218 240
R4542 VDD.n223 VDD.n222 240
R4543 VDD.n227 VDD.n226 240
R4544 VDD.n229 VDD.n150 240
R4545 VDD.n233 VDD.n129 240
R4546 VDD.n242 VDD.n127 240
R4547 VDD.n242 VDD.n122 240
R4548 VDD.n251 VDD.n122 240
R4549 VDD.n252 VDD.n251 240
R4550 VDD.n252 VDD.n66 240
R4551 VDD.n67 VDD.n66 240
R4552 VDD.n68 VDD.n67 240
R4553 VDD.n257 VDD.n68 240
R4554 VDD.n257 VDD.n73 240
R4555 VDD.n74 VDD.n73 240
R4556 VDD.n75 VDD.n74 240
R4557 VDD.n262 VDD.n75 240
R4558 VDD.n262 VDD.n80 240
R4559 VDD.n81 VDD.n80 240
R4560 VDD.n82 VDD.n81 240
R4561 VDD.n267 VDD.n82 240
R4562 VDD.n267 VDD.n87 240
R4563 VDD.n88 VDD.n87 240
R4564 VDD.n89 VDD.n88 240
R4565 VDD.n272 VDD.n89 240
R4566 VDD.n272 VDD.n94 240
R4567 VDD.n95 VDD.n94 240
R4568 VDD.n96 VDD.n95 240
R4569 VDD.n360 VDD.n98 240
R4570 VDD.n358 VDD.n357 240
R4571 VDD.n354 VDD.n353 240
R4572 VDD.n351 VDD.n102 240
R4573 VDD.n347 VDD.n345 240
R4574 VDD.n343 VDD.n104 240
R4575 VDD.n339 VDD.n337 240
R4576 VDD.n335 VDD.n106 240
R4577 VDD.n331 VDD.n329 240
R4578 VDD.n327 VDD.n108 240
R4579 VDD.n323 VDD.n321 240
R4580 VDD.n319 VDD.n110 240
R4581 VDD.n315 VDD.n313 240
R4582 VDD.n311 VDD.n112 240
R4583 VDD.n307 VDD.n305 240
R4584 VDD.n303 VDD.n114 240
R4585 VDD.n299 VDD.n297 240
R4586 VDD.n295 VDD.n116 240
R4587 VDD.n291 VDD.n289 240
R4588 VDD.n287 VDD.n118 240
R4589 VDD.n283 VDD.n281 240
R4590 VDD.n279 VDD.n120 240
R4591 VDD.n522 VDD.t86 231.595
R4592 VDD.n526 VDD.t49 231.595
R4593 VDD.n531 VDD.t60 231.595
R4594 VDD.n536 VDD.t95 231.595
R4595 VDD.n501 VDD.t88 231.595
R4596 VDD.n496 VDD.t54 231.595
R4597 VDD.n491 VDD.t45 231.595
R4598 VDD.t97 VDD.n486 231.595
R4599 VDD.n418 VDD.t75 231.595
R4600 VDD.n422 VDD.t66 231.595
R4601 VDD.n427 VDD.t63 231.595
R4602 VDD.n432 VDD.t42 231.595
R4603 VDD.n437 VDD.t57 231.595
R4604 VDD.n442 VDD.t69 231.595
R4605 VDD.n447 VDD.t52 231.595
R4606 VDD.n33 VDD.t81 231.595
R4607 VDD.n28 VDD.t92 231.595
R4608 VDD.n23 VDD.t83 231.595
R4609 VDD.n18 VDD.t77 231.595
R4610 VDD.n13 VDD.t90 231.595
R4611 VDD.n8 VDD.t72 231.595
R4612 VDD.n3 VDD.t79 231.595
R4613 VDD.n480 VDD.n478 204.214
R4614 VDD.n406 VDD.n404 204.214
R4615 VDD.n539 VDD.n538 203.03
R4616 VDD.n534 VDD.n533 203.03
R4617 VDD.n529 VDD.n528 203.03
R4618 VDD.n524 VDD.n523 203.03
R4619 VDD.n484 VDD.n483 203.03
R4620 VDD.n482 VDD.n481 203.03
R4621 VDD.n480 VDD.n479 203.03
R4622 VDD.n514 VDD.n513 203.03
R4623 VDD.n490 VDD.n488 203.03
R4624 VDD.n495 VDD.n493 203.03
R4625 VDD.n500 VDD.n498 203.03
R4626 VDD.n450 VDD.n449 203.03
R4627 VDD.n445 VDD.n444 203.03
R4628 VDD.n440 VDD.n439 203.03
R4629 VDD.n435 VDD.n434 203.03
R4630 VDD.n430 VDD.n429 203.03
R4631 VDD.n425 VDD.n424 203.03
R4632 VDD.n420 VDD.n419 203.03
R4633 VDD.n416 VDD.n415 203.03
R4634 VDD.n414 VDD.n413 203.03
R4635 VDD.n412 VDD.n411 203.03
R4636 VDD.n410 VDD.n409 203.03
R4637 VDD.n408 VDD.n407 203.03
R4638 VDD.n406 VDD.n405 203.03
R4639 VDD.n2 VDD.n1 203.03
R4640 VDD.n7 VDD.n5 203.03
R4641 VDD.n12 VDD.n10 203.03
R4642 VDD.n17 VDD.n15 203.03
R4643 VDD.n22 VDD.n20 203.03
R4644 VDD.n27 VDD.n25 203.03
R4645 VDD.n32 VDD.n30 203.03
R4646 VDD.n800 VDD.n799 185
R4647 VDD.n799 VDD.n798 185
R4648 VDD.n558 VDD.n556 185
R4649 VDD.n574 VDD.n573 185
R4650 VDD.n576 VDD.n575 185
R4651 VDD.n578 VDD.n577 185
R4652 VDD.n580 VDD.n579 185
R4653 VDD.n582 VDD.n581 185
R4654 VDD.n584 VDD.n583 185
R4655 VDD.n586 VDD.n585 185
R4656 VDD.n588 VDD.n587 185
R4657 VDD.n590 VDD.n589 185
R4658 VDD.n592 VDD.n591 185
R4659 VDD.n594 VDD.n593 185
R4660 VDD.n596 VDD.n595 185
R4661 VDD.n598 VDD.n597 185
R4662 VDD.n600 VDD.n599 185
R4663 VDD.n602 VDD.n601 185
R4664 VDD.n604 VDD.n603 185
R4665 VDD.n606 VDD.n605 185
R4666 VDD.n608 VDD.n607 185
R4667 VDD.n610 VDD.n609 185
R4668 VDD.n612 VDD.n611 185
R4669 VDD.n614 VDD.n613 185
R4670 VDD.n615 VDD.n571 185
R4671 VDD.n796 VDD.n795 185
R4672 VDD.n794 VDD.n572 185
R4673 VDD.n572 VDD.n559 185
R4674 VDD.n793 VDD.n792 185
R4675 VDD.n792 VDD.n791 185
R4676 VDD.n617 VDD.n616 185
R4677 VDD.n784 VDD.n617 185
R4678 VDD.n783 VDD.n782 185
R4679 VDD.n785 VDD.n783 185
R4680 VDD.n781 VDD.n622 185
R4681 VDD.n622 VDD.n621 185
R4682 VDD.n780 VDD.n779 185
R4683 VDD.n779 VDD.n778 185
R4684 VDD.n624 VDD.n623 185
R4685 VDD.n771 VDD.n624 185
R4686 VDD.n770 VDD.n769 185
R4687 VDD.n772 VDD.n770 185
R4688 VDD.n768 VDD.n629 185
R4689 VDD.n629 VDD.n628 185
R4690 VDD.n767 VDD.n766 185
R4691 VDD.n766 VDD.n765 185
R4692 VDD.n631 VDD.n630 185
R4693 VDD.n758 VDD.n631 185
R4694 VDD.n757 VDD.n756 185
R4695 VDD.n759 VDD.n757 185
R4696 VDD.n755 VDD.n636 185
R4697 VDD.n636 VDD.n635 185
R4698 VDD.n754 VDD.n753 185
R4699 VDD.n753 VDD.n752 185
R4700 VDD.n638 VDD.n637 185
R4701 VDD.n745 VDD.n638 185
R4702 VDD.n744 VDD.n743 185
R4703 VDD.n746 VDD.n744 185
R4704 VDD.n742 VDD.n643 185
R4705 VDD.n643 VDD.n642 185
R4706 VDD.n741 VDD.n740 185
R4707 VDD.n740 VDD.n739 185
R4708 VDD.n645 VDD.n644 185
R4709 VDD.n646 VDD.n645 185
R4710 VDD.n732 VDD.n731 185
R4711 VDD.n733 VDD.n732 185
R4712 VDD.n730 VDD.n651 185
R4713 VDD.n651 VDD.n650 185
R4714 VDD.n729 VDD.n728 185
R4715 VDD.n728 VDD.n727 185
R4716 VDD.n653 VDD.n652 185
R4717 VDD.n654 VDD.n653 185
R4718 VDD.n720 VDD.n719 185
R4719 VDD.n721 VDD.n720 185
R4720 VDD.n718 VDD.n659 185
R4721 VDD.n717 VDD.n716 185
R4722 VDD.n714 VDD.n660 185
R4723 VDD.n712 VDD.n711 185
R4724 VDD.n710 VDD.n661 185
R4725 VDD.n709 VDD.n708 185
R4726 VDD.n706 VDD.n662 185
R4727 VDD.n704 VDD.n703 185
R4728 VDD.n702 VDD.n663 185
R4729 VDD.n701 VDD.n700 185
R4730 VDD.n698 VDD.n664 185
R4731 VDD.n696 VDD.n695 185
R4732 VDD.n694 VDD.n665 185
R4733 VDD.n693 VDD.n692 185
R4734 VDD.n690 VDD.n666 185
R4735 VDD.n688 VDD.n687 185
R4736 VDD.n686 VDD.n667 185
R4737 VDD.n685 VDD.n684 185
R4738 VDD.n682 VDD.n668 185
R4739 VDD.n680 VDD.n679 185
R4740 VDD.n678 VDD.n669 185
R4741 VDD.n677 VDD.n676 185
R4742 VDD.n674 VDD.n670 185
R4743 VDD.n672 VDD.n671 185
R4744 VDD.n657 VDD.n656 185
R4745 VDD.n658 VDD.n657 185
R4746 VDD.n723 VDD.n722 185
R4747 VDD.n722 VDD.n721 185
R4748 VDD.n724 VDD.n655 185
R4749 VDD.n655 VDD.n654 185
R4750 VDD.n726 VDD.n725 185
R4751 VDD.n727 VDD.n726 185
R4752 VDD.n649 VDD.n648 185
R4753 VDD.n650 VDD.n649 185
R4754 VDD.n735 VDD.n734 185
R4755 VDD.n734 VDD.n733 185
R4756 VDD.n736 VDD.n647 185
R4757 VDD.n647 VDD.n646 185
R4758 VDD.n738 VDD.n737 185
R4759 VDD.n739 VDD.n738 185
R4760 VDD.n641 VDD.n640 185
R4761 VDD.n642 VDD.n641 185
R4762 VDD.n748 VDD.n747 185
R4763 VDD.n747 VDD.n746 185
R4764 VDD.n749 VDD.n639 185
R4765 VDD.n745 VDD.n639 185
R4766 VDD.n751 VDD.n750 185
R4767 VDD.n752 VDD.n751 185
R4768 VDD.n634 VDD.n633 185
R4769 VDD.n635 VDD.n634 185
R4770 VDD.n761 VDD.n760 185
R4771 VDD.n760 VDD.n759 185
R4772 VDD.n762 VDD.n632 185
R4773 VDD.n758 VDD.n632 185
R4774 VDD.n764 VDD.n763 185
R4775 VDD.n765 VDD.n764 185
R4776 VDD.n627 VDD.n626 185
R4777 VDD.n628 VDD.n627 185
R4778 VDD.n774 VDD.n773 185
R4779 VDD.n773 VDD.n772 185
R4780 VDD.n775 VDD.n625 185
R4781 VDD.n771 VDD.n625 185
R4782 VDD.n777 VDD.n776 185
R4783 VDD.n778 VDD.n777 185
R4784 VDD.n620 VDD.n619 185
R4785 VDD.n621 VDD.n620 185
R4786 VDD.n787 VDD.n786 185
R4787 VDD.n786 VDD.n785 185
R4788 VDD.n788 VDD.n618 185
R4789 VDD.n784 VDD.n618 185
R4790 VDD.n790 VDD.n789 185
R4791 VDD.n791 VDD.n790 185
R4792 VDD.n557 VDD.n555 185
R4793 VDD.n559 VDD.n557 185
R4794 VDD.n362 VDD.n98 185
R4795 VDD.n98 VDD.n97 185
R4796 VDD.n361 VDD.n360 185
R4797 VDD.n358 VDD.n99 185
R4798 VDD.n357 VDD.n356 185
R4799 VDD.n355 VDD.n354 185
R4800 VDD.n353 VDD.n101 185
R4801 VDD.n351 VDD.n350 185
R4802 VDD.n349 VDD.n102 185
R4803 VDD.n348 VDD.n347 185
R4804 VDD.n345 VDD.n103 185
R4805 VDD.n343 VDD.n342 185
R4806 VDD.n341 VDD.n104 185
R4807 VDD.n340 VDD.n339 185
R4808 VDD.n337 VDD.n105 185
R4809 VDD.n335 VDD.n334 185
R4810 VDD.n333 VDD.n106 185
R4811 VDD.n332 VDD.n331 185
R4812 VDD.n329 VDD.n107 185
R4813 VDD.n327 VDD.n326 185
R4814 VDD.n325 VDD.n108 185
R4815 VDD.n324 VDD.n323 185
R4816 VDD.n321 VDD.n109 185
R4817 VDD.n319 VDD.n318 185
R4818 VDD.n317 VDD.n110 185
R4819 VDD.n316 VDD.n315 185
R4820 VDD.n313 VDD.n111 185
R4821 VDD.n311 VDD.n310 185
R4822 VDD.n309 VDD.n112 185
R4823 VDD.n308 VDD.n307 185
R4824 VDD.n305 VDD.n113 185
R4825 VDD.n303 VDD.n302 185
R4826 VDD.n301 VDD.n114 185
R4827 VDD.n300 VDD.n299 185
R4828 VDD.n297 VDD.n115 185
R4829 VDD.n295 VDD.n294 185
R4830 VDD.n293 VDD.n116 185
R4831 VDD.n292 VDD.n291 185
R4832 VDD.n289 VDD.n117 185
R4833 VDD.n287 VDD.n286 185
R4834 VDD.n285 VDD.n118 185
R4835 VDD.n284 VDD.n283 185
R4836 VDD.n281 VDD.n119 185
R4837 VDD.n279 VDD.n278 185
R4838 VDD.n277 VDD.n120 185
R4839 VDD.n120 VDD.n97 185
R4840 VDD.n276 VDD.n96 185
R4841 VDD.n365 VDD.n96 185
R4842 VDD.n275 VDD.n95 185
R4843 VDD.n366 VDD.n95 185
R4844 VDD.n274 VDD.n94 185
R4845 VDD.n367 VDD.n94 185
R4846 VDD.n273 VDD.n272 185
R4847 VDD.n272 VDD.n90 185
R4848 VDD.n271 VDD.n89 185
R4849 VDD.n373 VDD.n89 185
R4850 VDD.n270 VDD.n88 185
R4851 VDD.n374 VDD.n88 185
R4852 VDD.n269 VDD.n87 185
R4853 VDD.n375 VDD.n87 185
R4854 VDD.n268 VDD.n267 185
R4855 VDD.n267 VDD.n83 185
R4856 VDD.n266 VDD.n82 185
R4857 VDD.n381 VDD.n82 185
R4858 VDD.n265 VDD.n81 185
R4859 VDD.n382 VDD.n81 185
R4860 VDD.n264 VDD.n80 185
R4861 VDD.n383 VDD.n80 185
R4862 VDD.n263 VDD.n262 185
R4863 VDD.n262 VDD.n76 185
R4864 VDD.n261 VDD.n75 185
R4865 VDD.n389 VDD.n75 185
R4866 VDD.n260 VDD.n74 185
R4867 VDD.n390 VDD.n74 185
R4868 VDD.n259 VDD.n73 185
R4869 VDD.n391 VDD.n73 185
R4870 VDD.n258 VDD.n257 185
R4871 VDD.n257 VDD.n69 185
R4872 VDD.n256 VDD.n68 185
R4873 VDD.n397 VDD.n68 185
R4874 VDD.n255 VDD.n67 185
R4875 VDD.n398 VDD.n67 185
R4876 VDD.n254 VDD.n66 185
R4877 VDD.n399 VDD.n66 185
R4878 VDD.n253 VDD.n252 185
R4879 VDD.n252 VDD.n65 185
R4880 VDD.n251 VDD.n121 185
R4881 VDD.n251 VDD.n250 185
R4882 VDD.n240 VDD.n122 185
R4883 VDD.n243 VDD.n122 185
R4884 VDD.n242 VDD.n241 185
R4885 VDD.n244 VDD.n242 185
R4886 VDD.n239 VDD.n127 185
R4887 VDD.n127 VDD.n126 185
R4888 VDD.n238 VDD.n237 185
R4889 VDD.n129 VDD.n128 185
R4890 VDD.n233 VDD.n232 185
R4891 VDD.n231 VDD.n150 185
R4892 VDD.n230 VDD.n229 185
R4893 VDD.n228 VDD.n227 185
R4894 VDD.n226 VDD.n225 185
R4895 VDD.n224 VDD.n223 185
R4896 VDD.n222 VDD.n221 185
R4897 VDD.n220 VDD.n219 185
R4898 VDD.n218 VDD.n217 185
R4899 VDD.n216 VDD.n215 185
R4900 VDD.n214 VDD.n213 185
R4901 VDD.n212 VDD.n211 185
R4902 VDD.n210 VDD.n209 185
R4903 VDD.n208 VDD.n207 185
R4904 VDD.n206 VDD.n205 185
R4905 VDD.n204 VDD.n203 185
R4906 VDD.n202 VDD.n201 185
R4907 VDD.n200 VDD.n199 185
R4908 VDD.n198 VDD.n197 185
R4909 VDD.n196 VDD.n195 185
R4910 VDD.n194 VDD.n193 185
R4911 VDD.n192 VDD.n191 185
R4912 VDD.n190 VDD.n189 185
R4913 VDD.n188 VDD.n187 185
R4914 VDD.n186 VDD.n185 185
R4915 VDD.n184 VDD.n183 185
R4916 VDD.n182 VDD.n181 185
R4917 VDD.n180 VDD.n179 185
R4918 VDD.n178 VDD.n177 185
R4919 VDD.n176 VDD.n175 185
R4920 VDD.n174 VDD.n173 185
R4921 VDD.n172 VDD.n171 185
R4922 VDD.n170 VDD.n169 185
R4923 VDD.n168 VDD.n167 185
R4924 VDD.n166 VDD.n165 185
R4925 VDD.n164 VDD.n163 185
R4926 VDD.n162 VDD.n161 185
R4927 VDD.n160 VDD.n159 185
R4928 VDD.n158 VDD.n157 185
R4929 VDD.n156 VDD.n155 185
R4930 VDD.n154 VDD.n153 185
R4931 VDD.n152 VDD.n151 185
R4932 VDD.n125 VDD.n124 185
R4933 VDD.n126 VDD.n125 185
R4934 VDD.n246 VDD.n245 185
R4935 VDD.n245 VDD.n244 185
R4936 VDD.n247 VDD.n123 185
R4937 VDD.n243 VDD.n123 185
R4938 VDD.n249 VDD.n248 185
R4939 VDD.n250 VDD.n249 185
R4940 VDD.n63 VDD.n61 185
R4941 VDD.n65 VDD.n63 185
R4942 VDD.n401 VDD.n400 185
R4943 VDD.n400 VDD.n399 185
R4944 VDD.n64 VDD.n62 185
R4945 VDD.n398 VDD.n64 185
R4946 VDD.n396 VDD.n395 185
R4947 VDD.n397 VDD.n396 185
R4948 VDD.n394 VDD.n70 185
R4949 VDD.n70 VDD.n69 185
R4950 VDD.n393 VDD.n392 185
R4951 VDD.n392 VDD.n391 185
R4952 VDD.n72 VDD.n71 185
R4953 VDD.n390 VDD.n72 185
R4954 VDD.n388 VDD.n387 185
R4955 VDD.n389 VDD.n388 185
R4956 VDD.n386 VDD.n77 185
R4957 VDD.n77 VDD.n76 185
R4958 VDD.n385 VDD.n384 185
R4959 VDD.n384 VDD.n383 185
R4960 VDD.n79 VDD.n78 185
R4961 VDD.n382 VDD.n79 185
R4962 VDD.n380 VDD.n379 185
R4963 VDD.n381 VDD.n380 185
R4964 VDD.n378 VDD.n84 185
R4965 VDD.n84 VDD.n83 185
R4966 VDD.n377 VDD.n376 185
R4967 VDD.n376 VDD.n375 185
R4968 VDD.n86 VDD.n85 185
R4969 VDD.n374 VDD.n86 185
R4970 VDD.n372 VDD.n371 185
R4971 VDD.n373 VDD.n372 185
R4972 VDD.n370 VDD.n91 185
R4973 VDD.n91 VDD.n90 185
R4974 VDD.n369 VDD.n368 185
R4975 VDD.n368 VDD.n367 185
R4976 VDD.n93 VDD.n92 185
R4977 VDD.n366 VDD.n93 185
R4978 VDD.n364 VDD.n363 185
R4979 VDD.n365 VDD.n364 185
R4980 VDD.n553 VDD.t84 113.526
R4981 VDD.t84 VDD.n552 113.526
R4982 VDD.n549 VDD.t46 113.526
R4983 VDD.t46 VDD.n548 113.526
R4984 VDD.n545 VDD.t58 113.526
R4985 VDD.t58 VDD.n544 113.526
R4986 VDD.n541 VDD.t93 113.526
R4987 VDD.t93 VDD.n540 113.526
R4988 VDD.n517 VDD.t96 113.526
R4989 VDD.t96 VDD.n516 113.526
R4990 VDD.n511 VDD.t43 113.526
R4991 VDD.t43 VDD.n510 113.526
R4992 VDD.n507 VDD.t53 113.526
R4993 VDD.t53 VDD.n506 113.526
R4994 VDD.n503 VDD.t87 113.526
R4995 VDD.t87 VDD.n502 113.526
R4996 VDD.n476 VDD.t73 113.526
R4997 VDD.t73 VDD.n475 113.526
R4998 VDD.n472 VDD.t64 113.526
R4999 VDD.t64 VDD.n471 113.526
R5000 VDD.n468 VDD.t61 113.526
R5001 VDD.t61 VDD.n467 113.526
R5002 VDD.n464 VDD.t39 113.526
R5003 VDD.t39 VDD.n463 113.526
R5004 VDD.n460 VDD.t55 113.526
R5005 VDD.t55 VDD.n459 113.526
R5006 VDD.n456 VDD.t67 113.526
R5007 VDD.t67 VDD.n455 113.526
R5008 VDD.n452 VDD.t50 113.526
R5009 VDD.t50 VDD.n451 113.526
R5010 VDD.n59 VDD.t78 113.526
R5011 VDD.t78 VDD.n58 113.526
R5012 VDD.n55 VDD.t70 113.526
R5013 VDD.t70 VDD.n54 113.526
R5014 VDD.n51 VDD.t89 113.526
R5015 VDD.t89 VDD.n50 113.526
R5016 VDD.n47 VDD.t76 113.526
R5017 VDD.t76 VDD.n46 113.526
R5018 VDD.n43 VDD.t82 113.526
R5019 VDD.t82 VDD.n42 113.526
R5020 VDD.n39 VDD.t91 113.526
R5021 VDD.t91 VDD.n38 113.526
R5022 VDD.n35 VDD.t80 113.526
R5023 VDD.t80 VDD.n34 113.526
R5024 VDD.n363 VDD.n362 80.9417
R5025 VDD.n277 VDD.n276 80.9417
R5026 VDD.n801 VDD.n800 78.6829
R5027 VDD.n795 VDD.n794 74.9181
R5028 VDD.n674 VDD.n673 72.7879
R5029 VDD.n675 VDD.n669 72.7879
R5030 VDD.n682 VDD.n681 72.7879
R5031 VDD.n683 VDD.n667 72.7879
R5032 VDD.n690 VDD.n689 72.7879
R5033 VDD.n691 VDD.n665 72.7879
R5034 VDD.n698 VDD.n697 72.7879
R5035 VDD.n699 VDD.n663 72.7879
R5036 VDD.n706 VDD.n705 72.7879
R5037 VDD.n707 VDD.n661 72.7879
R5038 VDD.n714 VDD.n713 72.7879
R5039 VDD.n715 VDD.n659 72.7879
R5040 VDD.n560 VDD.n558 72.7879
R5041 VDD.n575 VDD.n561 72.7879
R5042 VDD.n579 VDD.n562 72.7879
R5043 VDD.n583 VDD.n563 72.7879
R5044 VDD.n587 VDD.n564 72.7879
R5045 VDD.n591 VDD.n565 72.7879
R5046 VDD.n595 VDD.n566 72.7879
R5047 VDD.n599 VDD.n567 72.7879
R5048 VDD.n603 VDD.n568 72.7879
R5049 VDD.n607 VDD.n569 72.7879
R5050 VDD.n611 VDD.n570 72.7879
R5051 VDD.n797 VDD.n571 72.7879
R5052 VDD.n574 VDD.n560 72.7879
R5053 VDD.n578 VDD.n561 72.7879
R5054 VDD.n582 VDD.n562 72.7879
R5055 VDD.n586 VDD.n563 72.7879
R5056 VDD.n590 VDD.n564 72.7879
R5057 VDD.n594 VDD.n565 72.7879
R5058 VDD.n598 VDD.n566 72.7879
R5059 VDD.n602 VDD.n567 72.7879
R5060 VDD.n606 VDD.n568 72.7879
R5061 VDD.n610 VDD.n569 72.7879
R5062 VDD.n613 VDD.n570 72.7879
R5063 VDD.n797 VDD.n796 72.7879
R5064 VDD.n716 VDD.n715 72.7879
R5065 VDD.n713 VDD.n712 72.7879
R5066 VDD.n708 VDD.n707 72.7879
R5067 VDD.n705 VDD.n704 72.7879
R5068 VDD.n700 VDD.n699 72.7879
R5069 VDD.n697 VDD.n696 72.7879
R5070 VDD.n692 VDD.n691 72.7879
R5071 VDD.n689 VDD.n688 72.7879
R5072 VDD.n684 VDD.n683 72.7879
R5073 VDD.n681 VDD.n680 72.7879
R5074 VDD.n676 VDD.n675 72.7879
R5075 VDD.n673 VDD.n672 72.7879
R5076 VDD.n154 VDD.n130 72.7879
R5077 VDD.n158 VDD.n131 72.7879
R5078 VDD.n162 VDD.n132 72.7879
R5079 VDD.n166 VDD.n133 72.7879
R5080 VDD.n170 VDD.n134 72.7879
R5081 VDD.n174 VDD.n135 72.7879
R5082 VDD.n178 VDD.n136 72.7879
R5083 VDD.n182 VDD.n137 72.7879
R5084 VDD.n186 VDD.n138 72.7879
R5085 VDD.n190 VDD.n139 72.7879
R5086 VDD.n194 VDD.n140 72.7879
R5087 VDD.n198 VDD.n141 72.7879
R5088 VDD.n202 VDD.n142 72.7879
R5089 VDD.n206 VDD.n143 72.7879
R5090 VDD.n210 VDD.n144 72.7879
R5091 VDD.n214 VDD.n145 72.7879
R5092 VDD.n218 VDD.n146 72.7879
R5093 VDD.n222 VDD.n147 72.7879
R5094 VDD.n226 VDD.n148 72.7879
R5095 VDD.n229 VDD.n149 72.7879
R5096 VDD.n234 VDD.n233 72.7879
R5097 VDD.n237 VDD.n236 72.7879
R5098 VDD.n360 VDD.n359 72.7879
R5099 VDD.n357 VDD.n100 72.7879
R5100 VDD.n353 VDD.n352 72.7879
R5101 VDD.n346 VDD.n102 72.7879
R5102 VDD.n345 VDD.n344 72.7879
R5103 VDD.n338 VDD.n104 72.7879
R5104 VDD.n337 VDD.n336 72.7879
R5105 VDD.n330 VDD.n106 72.7879
R5106 VDD.n329 VDD.n328 72.7879
R5107 VDD.n322 VDD.n108 72.7879
R5108 VDD.n321 VDD.n320 72.7879
R5109 VDD.n314 VDD.n110 72.7879
R5110 VDD.n313 VDD.n312 72.7879
R5111 VDD.n306 VDD.n112 72.7879
R5112 VDD.n305 VDD.n304 72.7879
R5113 VDD.n298 VDD.n114 72.7879
R5114 VDD.n297 VDD.n296 72.7879
R5115 VDD.n290 VDD.n116 72.7879
R5116 VDD.n289 VDD.n288 72.7879
R5117 VDD.n282 VDD.n118 72.7879
R5118 VDD.n281 VDD.n280 72.7879
R5119 VDD.n359 VDD.n358 72.7879
R5120 VDD.n354 VDD.n100 72.7879
R5121 VDD.n352 VDD.n351 72.7879
R5122 VDD.n347 VDD.n346 72.7879
R5123 VDD.n344 VDD.n343 72.7879
R5124 VDD.n339 VDD.n338 72.7879
R5125 VDD.n336 VDD.n335 72.7879
R5126 VDD.n331 VDD.n330 72.7879
R5127 VDD.n328 VDD.n327 72.7879
R5128 VDD.n323 VDD.n322 72.7879
R5129 VDD.n320 VDD.n319 72.7879
R5130 VDD.n315 VDD.n314 72.7879
R5131 VDD.n312 VDD.n311 72.7879
R5132 VDD.n307 VDD.n306 72.7879
R5133 VDD.n304 VDD.n303 72.7879
R5134 VDD.n299 VDD.n298 72.7879
R5135 VDD.n296 VDD.n295 72.7879
R5136 VDD.n291 VDD.n290 72.7879
R5137 VDD.n288 VDD.n287 72.7879
R5138 VDD.n283 VDD.n282 72.7879
R5139 VDD.n280 VDD.n279 72.7879
R5140 VDD.n236 VDD.n129 72.7879
R5141 VDD.n234 VDD.n150 72.7879
R5142 VDD.n227 VDD.n149 72.7879
R5143 VDD.n223 VDD.n148 72.7879
R5144 VDD.n219 VDD.n147 72.7879
R5145 VDD.n215 VDD.n146 72.7879
R5146 VDD.n211 VDD.n145 72.7879
R5147 VDD.n207 VDD.n144 72.7879
R5148 VDD.n203 VDD.n143 72.7879
R5149 VDD.n199 VDD.n142 72.7879
R5150 VDD.n195 VDD.n141 72.7879
R5151 VDD.n191 VDD.n140 72.7879
R5152 VDD.n187 VDD.n139 72.7879
R5153 VDD.n183 VDD.n138 72.7879
R5154 VDD.n179 VDD.n137 72.7879
R5155 VDD.n175 VDD.n136 72.7879
R5156 VDD.n171 VDD.n135 72.7879
R5157 VDD.n167 VDD.n134 72.7879
R5158 VDD.n163 VDD.n133 72.7879
R5159 VDD.n159 VDD.n132 72.7879
R5160 VDD.n155 VDD.n131 72.7879
R5161 VDD.n151 VDD.n130 72.7879
R5162 VDD.n723 VDD.n656 70.4005
R5163 VDD.n239 VDD.n238 70.4005
R5164 VDD.n152 VDD.n124 70.4005
R5165 VDD.n719 VDD.n718 64.377
R5166 VDD.n798 VDD.n559 58.5822
R5167 VDD.n798 VDD.n560 56.1076
R5168 VDD.n798 VDD.n561 56.1076
R5169 VDD.n798 VDD.n562 56.1076
R5170 VDD.n798 VDD.n563 56.1076
R5171 VDD.n798 VDD.n564 56.1076
R5172 VDD.n798 VDD.n565 56.1076
R5173 VDD.n798 VDD.n566 56.1076
R5174 VDD.n798 VDD.n567 56.1076
R5175 VDD.n798 VDD.n568 56.1076
R5176 VDD.n798 VDD.n569 56.1076
R5177 VDD.n798 VDD.n570 56.1076
R5178 VDD.n798 VDD.n797 56.1076
R5179 VDD.n715 VDD.n658 56.1076
R5180 VDD.n713 VDD.n658 56.1076
R5181 VDD.n707 VDD.n658 56.1076
R5182 VDD.n705 VDD.n658 56.1076
R5183 VDD.n699 VDD.n658 56.1076
R5184 VDD.n697 VDD.n658 56.1076
R5185 VDD.n691 VDD.n658 56.1076
R5186 VDD.n689 VDD.n658 56.1076
R5187 VDD.n683 VDD.n658 56.1076
R5188 VDD.n681 VDD.n658 56.1076
R5189 VDD.n675 VDD.n658 56.1076
R5190 VDD.n673 VDD.n658 56.1076
R5191 VDD.n359 VDD.n97 56.1076
R5192 VDD.n100 VDD.n97 56.1076
R5193 VDD.n352 VDD.n97 56.1076
R5194 VDD.n346 VDD.n97 56.1076
R5195 VDD.n344 VDD.n97 56.1076
R5196 VDD.n338 VDD.n97 56.1076
R5197 VDD.n336 VDD.n97 56.1076
R5198 VDD.n330 VDD.n97 56.1076
R5199 VDD.n328 VDD.n97 56.1076
R5200 VDD.n322 VDD.n97 56.1076
R5201 VDD.n320 VDD.n97 56.1076
R5202 VDD.n314 VDD.n97 56.1076
R5203 VDD.n312 VDD.n97 56.1076
R5204 VDD.n306 VDD.n97 56.1076
R5205 VDD.n304 VDD.n97 56.1076
R5206 VDD.n298 VDD.n97 56.1076
R5207 VDD.n296 VDD.n97 56.1076
R5208 VDD.n290 VDD.n97 56.1076
R5209 VDD.n288 VDD.n97 56.1076
R5210 VDD.n282 VDD.n97 56.1076
R5211 VDD.n280 VDD.n97 56.1076
R5212 VDD.n236 VDD.n235 56.1076
R5213 VDD.n235 VDD.n234 56.1076
R5214 VDD.n235 VDD.n149 56.1076
R5215 VDD.n235 VDD.n148 56.1076
R5216 VDD.n235 VDD.n147 56.1076
R5217 VDD.n235 VDD.n146 56.1076
R5218 VDD.n235 VDD.n145 56.1076
R5219 VDD.n235 VDD.n144 56.1076
R5220 VDD.n235 VDD.n143 56.1076
R5221 VDD.n235 VDD.n142 56.1076
R5222 VDD.n235 VDD.n141 56.1076
R5223 VDD.n235 VDD.n140 56.1076
R5224 VDD.n235 VDD.n139 56.1076
R5225 VDD.n235 VDD.n138 56.1076
R5226 VDD.n235 VDD.n137 56.1076
R5227 VDD.n235 VDD.n136 56.1076
R5228 VDD.n235 VDD.n135 56.1076
R5229 VDD.n235 VDD.n134 56.1076
R5230 VDD.n235 VDD.n133 56.1076
R5231 VDD.n235 VDD.n132 56.1076
R5232 VDD.n235 VDD.n131 56.1076
R5233 VDD.n235 VDD.n130 56.1076
R5234 VDD.n721 VDD.n658 44.9131
R5235 VDD.n365 VDD.n97 35.0343
R5236 VDD.n721 VDD.n654 33.1968
R5237 VDD.n727 VDD.n654 33.1968
R5238 VDD.n733 VDD.n650 33.1968
R5239 VDD.n733 VDD.n646 33.1968
R5240 VDD.n739 VDD.n646 33.1968
R5241 VDD.n746 VDD.n642 33.1968
R5242 VDD.n746 VDD.n745 33.1968
R5243 VDD.n752 VDD.n635 33.1968
R5244 VDD.n759 VDD.n635 33.1968
R5245 VDD.n759 VDD.n758 33.1968
R5246 VDD.n765 VDD.n628 33.1968
R5247 VDD.n772 VDD.n628 33.1968
R5248 VDD.n772 VDD.n771 33.1968
R5249 VDD.n778 VDD.n621 33.1968
R5250 VDD.n785 VDD.n621 33.1968
R5251 VDD.n785 VDD.n784 33.1968
R5252 VDD.n791 VDD.n559 33.1968
R5253 VDD.t11 VDD.n642 32.7086
R5254 VDD.n538 VDD.t9 28.5655
R5255 VDD.n538 VDD.t94 28.5655
R5256 VDD.n533 VDD.t29 28.5655
R5257 VDD.n533 VDD.t59 28.5655
R5258 VDD.n528 VDD.t28 28.5655
R5259 VDD.n528 VDD.t48 28.5655
R5260 VDD.n523 VDD.t110 28.5655
R5261 VDD.n523 VDD.t85 28.5655
R5262 VDD.n483 VDD.t34 28.5655
R5263 VDD.n483 VDD.t1 28.5655
R5264 VDD.n481 VDD.t37 28.5655
R5265 VDD.n481 VDD.t4 28.5655
R5266 VDD.n479 VDD.t103 28.5655
R5267 VDD.n479 VDD.t22 28.5655
R5268 VDD.n478 VDD.t31 28.5655
R5269 VDD.n478 VDD.t10 28.5655
R5270 VDD.n513 VDD.t97 28.5655
R5271 VDD.n513 VDD.t106 28.5655
R5272 VDD.t45 VDD.n490 28.5655
R5273 VDD.n490 VDD.t21 28.5655
R5274 VDD.t54 VDD.n495 28.5655
R5275 VDD.n495 VDD.t109 28.5655
R5276 VDD.t88 VDD.n500 28.5655
R5277 VDD.n500 VDD.t12 28.5655
R5278 VDD.n449 VDD.t26 28.5655
R5279 VDD.n449 VDD.t51 28.5655
R5280 VDD.n444 VDD.t20 28.5655
R5281 VDD.n444 VDD.t68 28.5655
R5282 VDD.n439 VDD.t108 28.5655
R5283 VDD.n439 VDD.t56 28.5655
R5284 VDD.n434 VDD.t3 28.5655
R5285 VDD.n434 VDD.t41 28.5655
R5286 VDD.n429 VDD.t18 28.5655
R5287 VDD.n429 VDD.t62 28.5655
R5288 VDD.n424 VDD.t100 28.5655
R5289 VDD.n424 VDD.t65 28.5655
R5290 VDD.n419 VDD.t32 28.5655
R5291 VDD.n419 VDD.t74 28.5655
R5292 VDD.n415 VDD.t23 28.5655
R5293 VDD.n415 VDD.t35 28.5655
R5294 VDD.n413 VDD.t27 28.5655
R5295 VDD.n413 VDD.t24 28.5655
R5296 VDD.n411 VDD.t14 28.5655
R5297 VDD.n411 VDD.t107 28.5655
R5298 VDD.n409 VDD.t98 28.5655
R5299 VDD.n409 VDD.t7 28.5655
R5300 VDD.n407 VDD.t38 28.5655
R5301 VDD.n407 VDD.t6 28.5655
R5302 VDD.n405 VDD.t99 28.5655
R5303 VDD.n405 VDD.t102 28.5655
R5304 VDD.n404 VDD.t104 28.5655
R5305 VDD.n404 VDD.t36 28.5655
R5306 VDD.t79 VDD.n2 28.5655
R5307 VDD.n2 VDD.t17 28.5655
R5308 VDD.t72 VDD.n7 28.5655
R5309 VDD.n7 VDD.t33 28.5655
R5310 VDD.t90 VDD.n12 28.5655
R5311 VDD.n12 VDD.t16 28.5655
R5312 VDD.t77 VDD.n17 28.5655
R5313 VDD.n17 VDD.t101 28.5655
R5314 VDD.t83 VDD.n22 28.5655
R5315 VDD.n22 VDD.t105 28.5655
R5316 VDD.t92 VDD.n27 28.5655
R5317 VDD.n27 VDD.t19 28.5655
R5318 VDD.t81 VDD.n32 28.5655
R5319 VDD.n32 VDD.t25 28.5655
R5320 VDD.n235 VDD.n126 26.8597
R5321 VDD.n745 VDD.t30 26.8504
R5322 VDD.n791 VDD.t47 26.8504
R5323 VDD.t44 VDD.n650 25.8741
R5324 VDD.n800 VDD.n556 25.6005
R5325 VDD.n573 VDD.n556 25.6005
R5326 VDD.n576 VDD.n573 25.6005
R5327 VDD.n577 VDD.n576 25.6005
R5328 VDD.n580 VDD.n577 25.6005
R5329 VDD.n581 VDD.n580 25.6005
R5330 VDD.n584 VDD.n581 25.6005
R5331 VDD.n585 VDD.n584 25.6005
R5332 VDD.n588 VDD.n585 25.6005
R5333 VDD.n589 VDD.n588 25.6005
R5334 VDD.n592 VDD.n589 25.6005
R5335 VDD.n593 VDD.n592 25.6005
R5336 VDD.n596 VDD.n593 25.6005
R5337 VDD.n597 VDD.n596 25.6005
R5338 VDD.n600 VDD.n597 25.6005
R5339 VDD.n601 VDD.n600 25.6005
R5340 VDD.n604 VDD.n601 25.6005
R5341 VDD.n605 VDD.n604 25.6005
R5342 VDD.n608 VDD.n605 25.6005
R5343 VDD.n609 VDD.n608 25.6005
R5344 VDD.n612 VDD.n609 25.6005
R5345 VDD.n614 VDD.n612 25.6005
R5346 VDD.n615 VDD.n614 25.6005
R5347 VDD.n795 VDD.n615 25.6005
R5348 VDD.n719 VDD.n652 25.6005
R5349 VDD.n729 VDD.n652 25.6005
R5350 VDD.n730 VDD.n729 25.6005
R5351 VDD.n731 VDD.n730 25.6005
R5352 VDD.n731 VDD.n644 25.6005
R5353 VDD.n741 VDD.n644 25.6005
R5354 VDD.n742 VDD.n741 25.6005
R5355 VDD.n743 VDD.n742 25.6005
R5356 VDD.n743 VDD.n637 25.6005
R5357 VDD.n754 VDD.n637 25.6005
R5358 VDD.n755 VDD.n754 25.6005
R5359 VDD.n756 VDD.n755 25.6005
R5360 VDD.n756 VDD.n630 25.6005
R5361 VDD.n767 VDD.n630 25.6005
R5362 VDD.n768 VDD.n767 25.6005
R5363 VDD.n769 VDD.n768 25.6005
R5364 VDD.n769 VDD.n623 25.6005
R5365 VDD.n780 VDD.n623 25.6005
R5366 VDD.n781 VDD.n780 25.6005
R5367 VDD.n782 VDD.n781 25.6005
R5368 VDD.n782 VDD.n616 25.6005
R5369 VDD.n793 VDD.n616 25.6005
R5370 VDD.n794 VDD.n793 25.6005
R5371 VDD.n671 VDD.n656 25.6005
R5372 VDD.n671 VDD.n670 25.6005
R5373 VDD.n677 VDD.n670 25.6005
R5374 VDD.n678 VDD.n677 25.6005
R5375 VDD.n679 VDD.n678 25.6005
R5376 VDD.n679 VDD.n668 25.6005
R5377 VDD.n685 VDD.n668 25.6005
R5378 VDD.n686 VDD.n685 25.6005
R5379 VDD.n687 VDD.n686 25.6005
R5380 VDD.n687 VDD.n666 25.6005
R5381 VDD.n693 VDD.n666 25.6005
R5382 VDD.n694 VDD.n693 25.6005
R5383 VDD.n695 VDD.n694 25.6005
R5384 VDD.n695 VDD.n664 25.6005
R5385 VDD.n701 VDD.n664 25.6005
R5386 VDD.n702 VDD.n701 25.6005
R5387 VDD.n703 VDD.n702 25.6005
R5388 VDD.n703 VDD.n662 25.6005
R5389 VDD.n709 VDD.n662 25.6005
R5390 VDD.n710 VDD.n709 25.6005
R5391 VDD.n711 VDD.n710 25.6005
R5392 VDD.n711 VDD.n660 25.6005
R5393 VDD.n717 VDD.n660 25.6005
R5394 VDD.n718 VDD.n717 25.6005
R5395 VDD.n724 VDD.n723 25.6005
R5396 VDD.n725 VDD.n724 25.6005
R5397 VDD.n725 VDD.n648 25.6005
R5398 VDD.n735 VDD.n648 25.6005
R5399 VDD.n736 VDD.n735 25.6005
R5400 VDD.n737 VDD.n736 25.6005
R5401 VDD.n737 VDD.n640 25.6005
R5402 VDD.n748 VDD.n640 25.6005
R5403 VDD.n749 VDD.n748 25.6005
R5404 VDD.n750 VDD.n749 25.6005
R5405 VDD.n750 VDD.n633 25.6005
R5406 VDD.n761 VDD.n633 25.6005
R5407 VDD.n762 VDD.n761 25.6005
R5408 VDD.n763 VDD.n762 25.6005
R5409 VDD.n763 VDD.n626 25.6005
R5410 VDD.n774 VDD.n626 25.6005
R5411 VDD.n775 VDD.n774 25.6005
R5412 VDD.n776 VDD.n775 25.6005
R5413 VDD.n776 VDD.n619 25.6005
R5414 VDD.n787 VDD.n619 25.6005
R5415 VDD.n788 VDD.n787 25.6005
R5416 VDD.n789 VDD.n788 25.6005
R5417 VDD.n789 VDD.n555 25.6005
R5418 VDD.n362 VDD.n361 25.6005
R5419 VDD.n361 VDD.n99 25.6005
R5420 VDD.n356 VDD.n99 25.6005
R5421 VDD.n356 VDD.n355 25.6005
R5422 VDD.n355 VDD.n101 25.6005
R5423 VDD.n350 VDD.n101 25.6005
R5424 VDD.n350 VDD.n349 25.6005
R5425 VDD.n349 VDD.n348 25.6005
R5426 VDD.n348 VDD.n103 25.6005
R5427 VDD.n342 VDD.n103 25.6005
R5428 VDD.n342 VDD.n341 25.6005
R5429 VDD.n341 VDD.n340 25.6005
R5430 VDD.n340 VDD.n105 25.6005
R5431 VDD.n334 VDD.n105 25.6005
R5432 VDD.n334 VDD.n333 25.6005
R5433 VDD.n333 VDD.n332 25.6005
R5434 VDD.n332 VDD.n107 25.6005
R5435 VDD.n326 VDD.n107 25.6005
R5436 VDD.n326 VDD.n325 25.6005
R5437 VDD.n325 VDD.n324 25.6005
R5438 VDD.n324 VDD.n109 25.6005
R5439 VDD.n318 VDD.n109 25.6005
R5440 VDD.n318 VDD.n317 25.6005
R5441 VDD.n317 VDD.n316 25.6005
R5442 VDD.n316 VDD.n111 25.6005
R5443 VDD.n310 VDD.n111 25.6005
R5444 VDD.n310 VDD.n309 25.6005
R5445 VDD.n309 VDD.n308 25.6005
R5446 VDD.n308 VDD.n113 25.6005
R5447 VDD.n302 VDD.n113 25.6005
R5448 VDD.n302 VDD.n301 25.6005
R5449 VDD.n301 VDD.n300 25.6005
R5450 VDD.n300 VDD.n115 25.6005
R5451 VDD.n294 VDD.n115 25.6005
R5452 VDD.n294 VDD.n293 25.6005
R5453 VDD.n293 VDD.n292 25.6005
R5454 VDD.n292 VDD.n117 25.6005
R5455 VDD.n286 VDD.n117 25.6005
R5456 VDD.n286 VDD.n285 25.6005
R5457 VDD.n285 VDD.n284 25.6005
R5458 VDD.n284 VDD.n119 25.6005
R5459 VDD.n278 VDD.n119 25.6005
R5460 VDD.n278 VDD.n277 25.6005
R5461 VDD.n241 VDD.n239 25.6005
R5462 VDD.n241 VDD.n240 25.6005
R5463 VDD.n240 VDD.n121 25.6005
R5464 VDD.n253 VDD.n121 25.6005
R5465 VDD.n254 VDD.n253 25.6005
R5466 VDD.n255 VDD.n254 25.6005
R5467 VDD.n256 VDD.n255 25.6005
R5468 VDD.n258 VDD.n256 25.6005
R5469 VDD.n259 VDD.n258 25.6005
R5470 VDD.n260 VDD.n259 25.6005
R5471 VDD.n261 VDD.n260 25.6005
R5472 VDD.n263 VDD.n261 25.6005
R5473 VDD.n264 VDD.n263 25.6005
R5474 VDD.n265 VDD.n264 25.6005
R5475 VDD.n266 VDD.n265 25.6005
R5476 VDD.n268 VDD.n266 25.6005
R5477 VDD.n269 VDD.n268 25.6005
R5478 VDD.n270 VDD.n269 25.6005
R5479 VDD.n271 VDD.n270 25.6005
R5480 VDD.n273 VDD.n271 25.6005
R5481 VDD.n274 VDD.n273 25.6005
R5482 VDD.n275 VDD.n274 25.6005
R5483 VDD.n276 VDD.n275 25.6005
R5484 VDD.n153 VDD.n152 25.6005
R5485 VDD.n156 VDD.n153 25.6005
R5486 VDD.n157 VDD.n156 25.6005
R5487 VDD.n160 VDD.n157 25.6005
R5488 VDD.n161 VDD.n160 25.6005
R5489 VDD.n164 VDD.n161 25.6005
R5490 VDD.n165 VDD.n164 25.6005
R5491 VDD.n168 VDD.n165 25.6005
R5492 VDD.n169 VDD.n168 25.6005
R5493 VDD.n172 VDD.n169 25.6005
R5494 VDD.n173 VDD.n172 25.6005
R5495 VDD.n176 VDD.n173 25.6005
R5496 VDD.n177 VDD.n176 25.6005
R5497 VDD.n180 VDD.n177 25.6005
R5498 VDD.n181 VDD.n180 25.6005
R5499 VDD.n184 VDD.n181 25.6005
R5500 VDD.n185 VDD.n184 25.6005
R5501 VDD.n188 VDD.n185 25.6005
R5502 VDD.n189 VDD.n188 25.6005
R5503 VDD.n192 VDD.n189 25.6005
R5504 VDD.n193 VDD.n192 25.6005
R5505 VDD.n196 VDD.n193 25.6005
R5506 VDD.n197 VDD.n196 25.6005
R5507 VDD.n200 VDD.n197 25.6005
R5508 VDD.n201 VDD.n200 25.6005
R5509 VDD.n204 VDD.n201 25.6005
R5510 VDD.n205 VDD.n204 25.6005
R5511 VDD.n208 VDD.n205 25.6005
R5512 VDD.n209 VDD.n208 25.6005
R5513 VDD.n212 VDD.n209 25.6005
R5514 VDD.n213 VDD.n212 25.6005
R5515 VDD.n216 VDD.n213 25.6005
R5516 VDD.n217 VDD.n216 25.6005
R5517 VDD.n220 VDD.n217 25.6005
R5518 VDD.n221 VDD.n220 25.6005
R5519 VDD.n224 VDD.n221 25.6005
R5520 VDD.n225 VDD.n224 25.6005
R5521 VDD.n228 VDD.n225 25.6005
R5522 VDD.n230 VDD.n228 25.6005
R5523 VDD.n231 VDD.n230 25.6005
R5524 VDD.n232 VDD.n231 25.6005
R5525 VDD.n232 VDD.n128 25.6005
R5526 VDD.n238 VDD.n128 25.6005
R5527 VDD.n246 VDD.n124 25.6005
R5528 VDD.n247 VDD.n246 25.6005
R5529 VDD.n248 VDD.n247 25.6005
R5530 VDD.n248 VDD.n61 25.6005
R5531 VDD.n401 VDD.n62 25.6005
R5532 VDD.n395 VDD.n62 25.6005
R5533 VDD.n395 VDD.n394 25.6005
R5534 VDD.n394 VDD.n393 25.6005
R5535 VDD.n393 VDD.n71 25.6005
R5536 VDD.n387 VDD.n71 25.6005
R5537 VDD.n387 VDD.n386 25.6005
R5538 VDD.n386 VDD.n385 25.6005
R5539 VDD.n385 VDD.n78 25.6005
R5540 VDD.n379 VDD.n78 25.6005
R5541 VDD.n379 VDD.n378 25.6005
R5542 VDD.n378 VDD.n377 25.6005
R5543 VDD.n377 VDD.n85 25.6005
R5544 VDD.n371 VDD.n85 25.6005
R5545 VDD.n371 VDD.n370 25.6005
R5546 VDD.n370 VDD.n369 25.6005
R5547 VDD.n369 VDD.n92 25.6005
R5548 VDD.n363 VDD.n92 25.6005
R5549 VDD.n402 VDD.n401 22.5887
R5550 VDD.n805 VDD.n804 22.4706
R5551 VDD.n758 VDD.t0 20.0159
R5552 VDD.n778 VDD.t8 20.0159
R5553 VDD.n244 VDD.n126 19.853
R5554 VDD.n244 VDD.n243 19.853
R5555 VDD.n250 VDD.n65 19.853
R5556 VDD.n399 VDD.n65 19.853
R5557 VDD.n399 VDD.n398 19.853
R5558 VDD.n397 VDD.n69 19.853
R5559 VDD.n391 VDD.n69 19.853
R5560 VDD.n390 VDD.n389 19.853
R5561 VDD.n389 VDD.n76 19.853
R5562 VDD.n383 VDD.n76 19.853
R5563 VDD.n382 VDD.n381 19.853
R5564 VDD.n381 VDD.n83 19.853
R5565 VDD.n375 VDD.n83 19.853
R5566 VDD.n374 VDD.n373 19.853
R5567 VDD.n373 VDD.n90 19.853
R5568 VDD.n367 VDD.n90 19.853
R5569 VDD.n366 VDD.n365 19.853
R5570 VDD.t15 VDD.n397 19.561
R5571 VDD.n391 VDD.t13 16.0577
R5572 VDD.t40 VDD.n366 16.0577
R5573 VDD.n250 VDD.t71 15.4738
R5574 VDD.n765 VDD.t0 13.1814
R5575 VDD.n771 VDD.t8 13.1814
R5576 VDD.n383 VDD.t5 11.9704
R5577 VDD.t2 VDD.n374 11.9704
R5578 VDD VDD.n809 9.84561
R5579 VDD.n802 VDD.n801 9.3005
R5580 VDD.n403 VDD.n402 9.3005
R5581 VDD.t5 VDD.n382 7.88311
R5582 VDD.n375 VDD.t2 7.88311
R5583 VDD.n727 VDD.t44 7.32321
R5584 VDD.n752 VDD.t30 6.34685
R5585 VDD.n784 VDD.t47 6.34685
R5586 VDD.n243 VDD.t71 4.37973
R5587 VDD.t13 VDD.n390 3.79583
R5588 VDD.n367 VDD.t40 3.79583
R5589 VDD.n402 VDD.n61 3.01226
R5590 VDD.n801 VDD.n555 2.25932
R5591 VDD.n519 VDD.n518 1.45974
R5592 VDD.n520 VDD.n519 1.40267
R5593 VDD.n808 VDD.n807 1.40267
R5594 VDD.n807 VDD.n806 1.40267
R5595 VDD.n807 VDD.n416 1.40003
R5596 VDD.n804 VDD.n520 1.28854
R5597 VDD.n520 VDD.n484 1.26688
R5598 VDD.n803 VDD.n802 1.24507
R5599 VDD.n484 VDD.n482 1.18544
R5600 VDD.n482 VDD.n480 1.18544
R5601 VDD.n416 VDD.n414 1.18544
R5602 VDD.n414 VDD.n412 1.18544
R5603 VDD.n412 VDD.n410 1.18544
R5604 VDD.n410 VDD.n408 1.18544
R5605 VDD.n408 VDD.n406 1.18544
R5606 VDD.n805 VDD.n477 0.891804
R5607 VDD.n806 VDD.n417 0.891804
R5608 VDD.n809 VDD.n0 0.891804
R5609 VDD.n803 VDD.n521 0.758652
R5610 VDD.n519 VDD.n485 0.758652
R5611 VDD.n540 VDD.n539 0.734338
R5612 VDD.n540 VDD.n536 0.734338
R5613 VDD.n502 VDD.n501 0.734338
R5614 VDD.n502 VDD.n498 0.734338
R5615 VDD.n451 VDD.n450 0.734338
R5616 VDD.n451 VDD.n447 0.734338
R5617 VDD.n34 VDD.n33 0.734338
R5618 VDD.n34 VDD.n30 0.734338
R5619 VDD.n809 VDD.n808 0.701587
R5620 VDD.n806 VDD.n805 0.701587
R5621 VDD.n808 VDD.n403 0.67713
R5622 VDD.n739 VDD.t11 0.488681
R5623 VDD.n539 VDD.n537 0.38373
R5624 VDD.n542 VDD.n536 0.38373
R5625 VDD.n534 VDD.n532 0.38373
R5626 VDD.n546 VDD.n531 0.38373
R5627 VDD.n529 VDD.n527 0.38373
R5628 VDD.n550 VDD.n526 0.38373
R5629 VDD.n524 VDD.n521 0.38373
R5630 VDD.n554 VDD.n522 0.38373
R5631 VDD.n501 VDD.n499 0.38373
R5632 VDD.n504 VDD.n498 0.38373
R5633 VDD.n496 VDD.n494 0.38373
R5634 VDD.n508 VDD.n493 0.38373
R5635 VDD.n491 VDD.n489 0.38373
R5636 VDD.n512 VDD.n488 0.38373
R5637 VDD.n518 VDD.n486 0.38373
R5638 VDD.n514 VDD.n485 0.38373
R5639 VDD.n450 VDD.n448 0.38373
R5640 VDD.n453 VDD.n447 0.38373
R5641 VDD.n445 VDD.n443 0.38373
R5642 VDD.n457 VDD.n442 0.38373
R5643 VDD.n440 VDD.n438 0.38373
R5644 VDD.n461 VDD.n437 0.38373
R5645 VDD.n435 VDD.n433 0.38373
R5646 VDD.n465 VDD.n432 0.38373
R5647 VDD.n430 VDD.n428 0.38373
R5648 VDD.n469 VDD.n427 0.38373
R5649 VDD.n425 VDD.n423 0.38373
R5650 VDD.n473 VDD.n422 0.38373
R5651 VDD.n420 VDD.n417 0.38373
R5652 VDD.n477 VDD.n418 0.38373
R5653 VDD.n33 VDD.n31 0.38373
R5654 VDD.n36 VDD.n30 0.38373
R5655 VDD.n28 VDD.n26 0.38373
R5656 VDD.n40 VDD.n25 0.38373
R5657 VDD.n23 VDD.n21 0.38373
R5658 VDD.n44 VDD.n20 0.38373
R5659 VDD.n18 VDD.n16 0.38373
R5660 VDD.n48 VDD.n15 0.38373
R5661 VDD.n13 VDD.n11 0.38373
R5662 VDD.n52 VDD.n10 0.38373
R5663 VDD.n8 VDD.n6 0.38373
R5664 VDD.n56 VDD.n5 0.38373
R5665 VDD.n3 VDD.n0 0.38373
R5666 VDD.n60 VDD.n1 0.38373
R5667 VDD.n535 VDD.n534 0.383729
R5668 VDD.n543 VDD.n531 0.383729
R5669 VDD.n530 VDD.n529 0.383729
R5670 VDD.n547 VDD.n526 0.383729
R5671 VDD.n525 VDD.n524 0.383729
R5672 VDD.n551 VDD.n522 0.383729
R5673 VDD.n497 VDD.n496 0.383729
R5674 VDD.n505 VDD.n493 0.383729
R5675 VDD.n492 VDD.n491 0.383729
R5676 VDD.n509 VDD.n488 0.383729
R5677 VDD.n487 VDD.n486 0.383729
R5678 VDD.n515 VDD.n514 0.383729
R5679 VDD.n446 VDD.n445 0.383729
R5680 VDD.n454 VDD.n442 0.383729
R5681 VDD.n441 VDD.n440 0.383729
R5682 VDD.n458 VDD.n437 0.383729
R5683 VDD.n436 VDD.n435 0.383729
R5684 VDD.n462 VDD.n432 0.383729
R5685 VDD.n431 VDD.n430 0.383729
R5686 VDD.n466 VDD.n427 0.383729
R5687 VDD.n426 VDD.n425 0.383729
R5688 VDD.n470 VDD.n422 0.383729
R5689 VDD.n421 VDD.n420 0.383729
R5690 VDD.n474 VDD.n418 0.383729
R5691 VDD.n29 VDD.n28 0.383729
R5692 VDD.n37 VDD.n25 0.383729
R5693 VDD.n24 VDD.n23 0.383729
R5694 VDD.n41 VDD.n20 0.383729
R5695 VDD.n19 VDD.n18 0.383729
R5696 VDD.n45 VDD.n15 0.383729
R5697 VDD.n14 VDD.n13 0.383729
R5698 VDD.n49 VDD.n10 0.383729
R5699 VDD.n9 VDD.n8 0.383729
R5700 VDD.n53 VDD.n5 0.383729
R5701 VDD.n4 VDD.n3 0.383729
R5702 VDD.n57 VDD.n1 0.383729
R5703 VDD.n541 VDD.n537 0.351109
R5704 VDD.n542 VDD.n541 0.351109
R5705 VDD.n544 VDD.n535 0.351109
R5706 VDD.n544 VDD.n543 0.351109
R5707 VDD.n545 VDD.n532 0.351109
R5708 VDD.n546 VDD.n545 0.351109
R5709 VDD.n548 VDD.n530 0.351109
R5710 VDD.n548 VDD.n547 0.351109
R5711 VDD.n549 VDD.n527 0.351109
R5712 VDD.n550 VDD.n549 0.351109
R5713 VDD.n552 VDD.n525 0.351109
R5714 VDD.n552 VDD.n551 0.351109
R5715 VDD.n553 VDD.n521 0.351109
R5716 VDD.n554 VDD.n553 0.351109
R5717 VDD.n503 VDD.n499 0.351109
R5718 VDD.n504 VDD.n503 0.351109
R5719 VDD.n506 VDD.n497 0.351109
R5720 VDD.n506 VDD.n505 0.351109
R5721 VDD.n507 VDD.n494 0.351109
R5722 VDD.n508 VDD.n507 0.351109
R5723 VDD.n510 VDD.n492 0.351109
R5724 VDD.n510 VDD.n509 0.351109
R5725 VDD.n511 VDD.n489 0.351109
R5726 VDD.n512 VDD.n511 0.351109
R5727 VDD.n516 VDD.n487 0.351109
R5728 VDD.n516 VDD.n515 0.351109
R5729 VDD.n518 VDD.n517 0.351109
R5730 VDD.n517 VDD.n485 0.351109
R5731 VDD.n452 VDD.n448 0.351109
R5732 VDD.n453 VDD.n452 0.351109
R5733 VDD.n455 VDD.n446 0.351109
R5734 VDD.n455 VDD.n454 0.351109
R5735 VDD.n456 VDD.n443 0.351109
R5736 VDD.n457 VDD.n456 0.351109
R5737 VDD.n459 VDD.n441 0.351109
R5738 VDD.n459 VDD.n458 0.351109
R5739 VDD.n460 VDD.n438 0.351109
R5740 VDD.n461 VDD.n460 0.351109
R5741 VDD.n463 VDD.n436 0.351109
R5742 VDD.n463 VDD.n462 0.351109
R5743 VDD.n464 VDD.n433 0.351109
R5744 VDD.n465 VDD.n464 0.351109
R5745 VDD.n467 VDD.n431 0.351109
R5746 VDD.n467 VDD.n466 0.351109
R5747 VDD.n468 VDD.n428 0.351109
R5748 VDD.n469 VDD.n468 0.351109
R5749 VDD.n471 VDD.n426 0.351109
R5750 VDD.n471 VDD.n470 0.351109
R5751 VDD.n472 VDD.n423 0.351109
R5752 VDD.n473 VDD.n472 0.351109
R5753 VDD.n475 VDD.n421 0.351109
R5754 VDD.n475 VDD.n474 0.351109
R5755 VDD.n476 VDD.n417 0.351109
R5756 VDD.n477 VDD.n476 0.351109
R5757 VDD.n35 VDD.n31 0.351109
R5758 VDD.n36 VDD.n35 0.351109
R5759 VDD.n38 VDD.n29 0.351109
R5760 VDD.n38 VDD.n37 0.351109
R5761 VDD.n39 VDD.n26 0.351109
R5762 VDD.n40 VDD.n39 0.351109
R5763 VDD.n42 VDD.n24 0.351109
R5764 VDD.n42 VDD.n41 0.351109
R5765 VDD.n43 VDD.n21 0.351109
R5766 VDD.n44 VDD.n43 0.351109
R5767 VDD.n46 VDD.n19 0.351109
R5768 VDD.n46 VDD.n45 0.351109
R5769 VDD.n47 VDD.n16 0.351109
R5770 VDD.n48 VDD.n47 0.351109
R5771 VDD.n50 VDD.n14 0.351109
R5772 VDD.n50 VDD.n49 0.351109
R5773 VDD.n51 VDD.n11 0.351109
R5774 VDD.n52 VDD.n51 0.351109
R5775 VDD.n54 VDD.n9 0.351109
R5776 VDD.n54 VDD.n53 0.351109
R5777 VDD.n55 VDD.n6 0.351109
R5778 VDD.n56 VDD.n55 0.351109
R5779 VDD.n58 VDD.n4 0.351109
R5780 VDD.n58 VDD.n57 0.351109
R5781 VDD.n59 VDD.n0 0.351109
R5782 VDD.n60 VDD.n59 0.351109
R5783 VDD.n398 VDD.t15 0.292448
R5784 VDD.n802 VDD.n554 0.215174
R5785 VDD.n403 VDD.n60 0.215174
R5786 VDD.n543 VDD.n542 0.168978
R5787 VDD.n537 VDD.n535 0.168978
R5788 VDD.n547 VDD.n546 0.168978
R5789 VDD.n532 VDD.n530 0.168978
R5790 VDD.n551 VDD.n550 0.168978
R5791 VDD.n527 VDD.n525 0.168978
R5792 VDD.n505 VDD.n504 0.168978
R5793 VDD.n499 VDD.n497 0.168978
R5794 VDD.n509 VDD.n508 0.168978
R5795 VDD.n494 VDD.n492 0.168978
R5796 VDD.n515 VDD.n512 0.168978
R5797 VDD.n489 VDD.n487 0.168978
R5798 VDD.n454 VDD.n453 0.168978
R5799 VDD.n448 VDD.n446 0.168978
R5800 VDD.n458 VDD.n457 0.168978
R5801 VDD.n443 VDD.n441 0.168978
R5802 VDD.n462 VDD.n461 0.168978
R5803 VDD.n438 VDD.n436 0.168978
R5804 VDD.n466 VDD.n465 0.168978
R5805 VDD.n433 VDD.n431 0.168978
R5806 VDD.n470 VDD.n469 0.168978
R5807 VDD.n428 VDD.n426 0.168978
R5808 VDD.n474 VDD.n473 0.168978
R5809 VDD.n423 VDD.n421 0.168978
R5810 VDD.n37 VDD.n36 0.168978
R5811 VDD.n31 VDD.n29 0.168978
R5812 VDD.n41 VDD.n40 0.168978
R5813 VDD.n26 VDD.n24 0.168978
R5814 VDD.n45 VDD.n44 0.168978
R5815 VDD.n21 VDD.n19 0.168978
R5816 VDD.n49 VDD.n48 0.168978
R5817 VDD.n16 VDD.n14 0.168978
R5818 VDD.n53 VDD.n52 0.168978
R5819 VDD.n11 VDD.n9 0.168978
R5820 VDD.n57 VDD.n56 0.168978
R5821 VDD.n6 VDD.n4 0.168978
R5822 VDD.n804 VDD.n803 0.11463
R5823 IBIAS.n9 IBIAS.t42 117.266
R5824 IBIAS.n14 IBIAS.t20 117.266
R5825 IBIAS.n20 IBIAS.t46 117.266
R5826 IBIAS.n26 IBIAS.t40 117.266
R5827 IBIAS.n32 IBIAS.t74 117.266
R5828 IBIAS.n38 IBIAS.t70 117.266
R5829 IBIAS.n44 IBIAS.t108 117.266
R5830 IBIAS.n50 IBIAS.t73 117.266
R5831 IBIAS.n56 IBIAS.t109 117.266
R5832 IBIAS.n62 IBIAS.t34 117.266
R5833 IBIAS.n93 IBIAS.t27 117.266
R5834 IBIAS.n90 IBIAS.t80 117.266
R5835 IBIAS.n87 IBIAS.t53 117.266
R5836 IBIAS.n84 IBIAS.t81 117.266
R5837 IBIAS.n81 IBIAS.t52 117.266
R5838 IBIAS.n78 IBIAS.t15 117.266
R5839 IBIAS.n75 IBIAS.t86 117.266
R5840 IBIAS.n68 IBIAS.t60 117.266
R5841 IBIAS.n5 IBIAS.t0 116.647
R5842 IBIAS.n6 IBIAS.t2 116.647
R5843 IBIAS.n1 IBIAS.t4 116.647
R5844 IBIAS.n2 IBIAS.t6 116.647
R5845 IBIAS.n74 IBIAS.t59 116.647
R5846 IBIAS.n73 IBIAS.t14 116.647
R5847 IBIAS.n72 IBIAS.t13 116.647
R5848 IBIAS.n71 IBIAS.t10 116.647
R5849 IBIAS.n70 IBIAS.t107 116.647
R5850 IBIAS.n69 IBIAS.t36 116.647
R5851 IBIAS.n68 IBIAS.t61 116.647
R5852 IBIAS.n13 IBIAS.t38 116.647
R5853 IBIAS.n12 IBIAS.t16 116.647
R5854 IBIAS.n11 IBIAS.t19 116.647
R5855 IBIAS.n10 IBIAS.t102 116.647
R5856 IBIAS.n9 IBIAS.t69 116.647
R5857 IBIAS.n18 IBIAS.t89 116.647
R5858 IBIAS.n17 IBIAS.t64 116.647
R5859 IBIAS.n16 IBIAS.t66 116.647
R5860 IBIAS.n15 IBIAS.t58 116.647
R5861 IBIAS.n14 IBIAS.t21 116.647
R5862 IBIAS.n24 IBIAS.t35 116.647
R5863 IBIAS.n23 IBIAS.t37 116.647
R5864 IBIAS.n22 IBIAS.t39 116.647
R5865 IBIAS.n21 IBIAS.t17 116.647
R5866 IBIAS.n20 IBIAS.t72 116.647
R5867 IBIAS.n30 IBIAS.t18 116.647
R5868 IBIAS.n29 IBIAS.t90 116.647
R5869 IBIAS.n28 IBIAS.t91 116.647
R5870 IBIAS.n27 IBIAS.t83 116.647
R5871 IBIAS.n26 IBIAS.t43 116.647
R5872 IBIAS.n36 IBIAS.t62 116.647
R5873 IBIAS.n35 IBIAS.t63 116.647
R5874 IBIAS.n34 IBIAS.t65 116.647
R5875 IBIAS.n33 IBIAS.t44 116.647
R5876 IBIAS.n32 IBIAS.t104 116.647
R5877 IBIAS.n42 IBIAS.t47 116.647
R5878 IBIAS.n41 IBIAS.t22 116.647
R5879 IBIAS.n40 IBIAS.t25 116.647
R5880 IBIAS.n39 IBIAS.t11 116.647
R5881 IBIAS.n38 IBIAS.t75 116.647
R5882 IBIAS.n48 IBIAS.t93 116.647
R5883 IBIAS.n47 IBIAS.t96 116.647
R5884 IBIAS.n46 IBIAS.t98 116.647
R5885 IBIAS.n45 IBIAS.t76 116.647
R5886 IBIAS.n44 IBIAS.t32 116.647
R5887 IBIAS.n54 IBIAS.t48 116.647
R5888 IBIAS.n53 IBIAS.t24 116.647
R5889 IBIAS.n52 IBIAS.t26 116.647
R5890 IBIAS.n51 IBIAS.t12 116.647
R5891 IBIAS.n50 IBIAS.t79 116.647
R5892 IBIAS.n60 IBIAS.t94 116.647
R5893 IBIAS.n59 IBIAS.t97 116.647
R5894 IBIAS.n58 IBIAS.t99 116.647
R5895 IBIAS.n57 IBIAS.t77 116.647
R5896 IBIAS.n56 IBIAS.t33 116.647
R5897 IBIAS.n66 IBIAS.t68 116.647
R5898 IBIAS.n65 IBIAS.t50 116.647
R5899 IBIAS.n64 IBIAS.t67 116.647
R5900 IBIAS.n63 IBIAS.t49 116.647
R5901 IBIAS.n62 IBIAS.t51 116.647
R5902 IBIAS.n99 IBIAS.t23 116.647
R5903 IBIAS.n98 IBIAS.t84 116.647
R5904 IBIAS.n97 IBIAS.t82 116.647
R5905 IBIAS.n96 IBIAS.t78 116.647
R5906 IBIAS.n95 IBIAS.t71 116.647
R5907 IBIAS.n94 IBIAS.t106 116.647
R5908 IBIAS.n93 IBIAS.t28 116.647
R5909 IBIAS.n92 IBIAS.t92 116.647
R5910 IBIAS.n91 IBIAS.t54 116.647
R5911 IBIAS.n90 IBIAS.t41 116.647
R5912 IBIAS.n89 IBIAS.t103 116.647
R5913 IBIAS.n88 IBIAS.t100 116.647
R5914 IBIAS.n87 IBIAS.t56 116.647
R5915 IBIAS.n86 IBIAS.t95 116.647
R5916 IBIAS.n85 IBIAS.t55 116.647
R5917 IBIAS.n84 IBIAS.t45 116.647
R5918 IBIAS.n83 IBIAS.t105 116.647
R5919 IBIAS.n82 IBIAS.t101 116.647
R5920 IBIAS.n81 IBIAS.t57 116.647
R5921 IBIAS.n80 IBIAS.t29 116.647
R5922 IBIAS.n79 IBIAS.t88 116.647
R5923 IBIAS.n78 IBIAS.t85 116.647
R5924 IBIAS.n77 IBIAS.t31 116.647
R5925 IBIAS.n76 IBIAS.t30 116.647
R5926 IBIAS.n75 IBIAS.t87 116.647
R5927 IBIAS.n1 IBIAS.n0 72.4405
R5928 IBIAS.n4 IBIAS.n3 72.2205
R5929 IBIAS.n8 IBIAS.n7 72.2205
R5930 IBIAS.n108 IBIAS.n107 19.6468
R5931 IBIAS.n0 IBIAS.t5 17.4005
R5932 IBIAS.n0 IBIAS.t8 17.4005
R5933 IBIAS.n3 IBIAS.t1 17.4005
R5934 IBIAS.n3 IBIAS.t7 17.4005
R5935 IBIAS.n7 IBIAS.t9 17.4005
R5936 IBIAS.n7 IBIAS.t3 17.4005
R5937 IBIAS.n107 IBIAS.n67 15.3043
R5938 IBIAS.n19 IBIAS.n13 6.03305
R5939 IBIAS IBIAS.n108 4.11588
R5940 IBIAS.n19 IBIAS.n18 3.91286
R5941 IBIAS.n31 IBIAS.n30 3.91286
R5942 IBIAS.n43 IBIAS.n42 3.91286
R5943 IBIAS.n55 IBIAS.n54 3.91286
R5944 IBIAS.n67 IBIAS.n66 3.91286
R5945 IBIAS.n101 IBIAS.n89 3.88358
R5946 IBIAS.n103 IBIAS.n83 3.88358
R5947 IBIAS.n105 IBIAS.n77 3.88358
R5948 IBIAS.n100 IBIAS.n99 3.58059
R5949 IBIAS.n25 IBIAS.n24 2.67247
R5950 IBIAS.n37 IBIAS.n36 2.67247
R5951 IBIAS.n49 IBIAS.n48 2.67247
R5952 IBIAS.n61 IBIAS.n60 2.67247
R5953 IBIAS.n106 IBIAS.n74 2.64347
R5954 IBIAS.n100 IBIAS.n92 2.6432
R5955 IBIAS.n102 IBIAS.n86 2.6432
R5956 IBIAS.n104 IBIAS.n80 2.6432
R5957 IBIAS.n15 IBIAS.n14 1.85887
R5958 IBIAS.n17 IBIAS.n16 1.85887
R5959 IBIAS.n21 IBIAS.n20 1.85887
R5960 IBIAS.n23 IBIAS.n22 1.85887
R5961 IBIAS.n27 IBIAS.n26 1.85887
R5962 IBIAS.n29 IBIAS.n28 1.85887
R5963 IBIAS.n33 IBIAS.n32 1.85887
R5964 IBIAS.n35 IBIAS.n34 1.85887
R5965 IBIAS.n39 IBIAS.n38 1.85887
R5966 IBIAS.n41 IBIAS.n40 1.85887
R5967 IBIAS.n45 IBIAS.n44 1.85887
R5968 IBIAS.n47 IBIAS.n46 1.85887
R5969 IBIAS.n51 IBIAS.n50 1.85887
R5970 IBIAS.n53 IBIAS.n52 1.85887
R5971 IBIAS.n57 IBIAS.n56 1.85887
R5972 IBIAS.n59 IBIAS.n58 1.85887
R5973 IBIAS.n91 IBIAS.n90 1.85887
R5974 IBIAS.n88 IBIAS.n87 1.85887
R5975 IBIAS.n85 IBIAS.n84 1.85887
R5976 IBIAS.n82 IBIAS.n81 1.85887
R5977 IBIAS.n79 IBIAS.n78 1.85887
R5978 IBIAS.n76 IBIAS.n75 1.85887
R5979 IBIAS.n107 IBIAS.n106 1.83961
R5980 IBIAS.n108 IBIAS.n8 1.42358
R5981 IBIAS.n101 IBIAS.n100 0.938028
R5982 IBIAS.n102 IBIAS.n101 0.938028
R5983 IBIAS.n103 IBIAS.n102 0.938028
R5984 IBIAS.n104 IBIAS.n103 0.938028
R5985 IBIAS.n105 IBIAS.n104 0.938028
R5986 IBIAS.n106 IBIAS.n105 0.937009
R5987 IBIAS.n25 IBIAS.n19 0.880308
R5988 IBIAS.n31 IBIAS.n25 0.880308
R5989 IBIAS.n37 IBIAS.n31 0.880308
R5990 IBIAS.n43 IBIAS.n37 0.880308
R5991 IBIAS.n49 IBIAS.n43 0.880308
R5992 IBIAS.n55 IBIAS.n49 0.880308
R5993 IBIAS.n61 IBIAS.n55 0.880308
R5994 IBIAS.n67 IBIAS.n61 0.880308
R5995 IBIAS.n2 IBIAS.n1 0.618487
R5996 IBIAS.n6 IBIAS.n5 0.618487
R5997 IBIAS.n10 IBIAS.n9 0.618487
R5998 IBIAS.n11 IBIAS.n10 0.618487
R5999 IBIAS.n12 IBIAS.n11 0.618487
R6000 IBIAS.n13 IBIAS.n12 0.618487
R6001 IBIAS.n16 IBIAS.n15 0.618487
R6002 IBIAS.n18 IBIAS.n17 0.618487
R6003 IBIAS.n22 IBIAS.n21 0.618487
R6004 IBIAS.n24 IBIAS.n23 0.618487
R6005 IBIAS.n28 IBIAS.n27 0.618487
R6006 IBIAS.n30 IBIAS.n29 0.618487
R6007 IBIAS.n34 IBIAS.n33 0.618487
R6008 IBIAS.n36 IBIAS.n35 0.618487
R6009 IBIAS.n40 IBIAS.n39 0.618487
R6010 IBIAS.n42 IBIAS.n41 0.618487
R6011 IBIAS.n46 IBIAS.n45 0.618487
R6012 IBIAS.n48 IBIAS.n47 0.618487
R6013 IBIAS.n52 IBIAS.n51 0.618487
R6014 IBIAS.n54 IBIAS.n53 0.618487
R6015 IBIAS.n58 IBIAS.n57 0.618487
R6016 IBIAS.n60 IBIAS.n59 0.618487
R6017 IBIAS.n63 IBIAS.n62 0.618487
R6018 IBIAS.n64 IBIAS.n63 0.618487
R6019 IBIAS.n65 IBIAS.n64 0.618487
R6020 IBIAS.n66 IBIAS.n65 0.618487
R6021 IBIAS.n94 IBIAS.n93 0.618487
R6022 IBIAS.n95 IBIAS.n94 0.618487
R6023 IBIAS.n96 IBIAS.n95 0.618487
R6024 IBIAS.n97 IBIAS.n96 0.618487
R6025 IBIAS.n98 IBIAS.n97 0.618487
R6026 IBIAS.n99 IBIAS.n98 0.618487
R6027 IBIAS.n92 IBIAS.n91 0.618487
R6028 IBIAS.n89 IBIAS.n88 0.618487
R6029 IBIAS.n86 IBIAS.n85 0.618487
R6030 IBIAS.n83 IBIAS.n82 0.618487
R6031 IBIAS.n80 IBIAS.n79 0.618487
R6032 IBIAS.n77 IBIAS.n76 0.618487
R6033 IBIAS.n69 IBIAS.n68 0.618487
R6034 IBIAS.n70 IBIAS.n69 0.618487
R6035 IBIAS.n71 IBIAS.n70 0.618487
R6036 IBIAS.n72 IBIAS.n71 0.618487
R6037 IBIAS.n73 IBIAS.n72 0.618487
R6038 IBIAS.n74 IBIAS.n73 0.618487
R6039 IBIAS.n4 IBIAS.n2 0.220551
R6040 IBIAS.n8 IBIAS.n6 0.220551
R6041 IBIAS.n5 IBIAS.n4 0.220551
R6042 a_3329_8823.n77 a_3329_8823.n76 76.1488
R6043 a_3329_8823.n5 a_3329_8823.n3 76.1487
R6044 a_3329_8823.n2 a_3329_8823.n0 76.1487
R6045 a_3329_8823.n57 a_3329_8823.n55 76.1487
R6046 a_3329_8823.n60 a_3329_8823.n58 76.1487
R6047 a_3329_8823.n63 a_3329_8823.n61 76.1487
R6048 a_3329_8823.n8 a_3329_8823.n6 75.8119
R6049 a_3329_8823.n66 a_3329_8823.n64 75.8119
R6050 a_3329_8823.n76 a_3329_8823.n75 75.4751
R6051 a_3329_8823.n12 a_3329_8823.n11 75.4751
R6052 a_3329_8823.n10 a_3329_8823.n9 75.4751
R6053 a_3329_8823.n8 a_3329_8823.n7 75.4751
R6054 a_3329_8823.n5 a_3329_8823.n4 75.4751
R6055 a_3329_8823.n2 a_3329_8823.n1 75.4751
R6056 a_3329_8823.n57 a_3329_8823.n56 75.4751
R6057 a_3329_8823.n60 a_3329_8823.n59 75.4751
R6058 a_3329_8823.n63 a_3329_8823.n62 75.4751
R6059 a_3329_8823.n70 a_3329_8823.n69 75.4751
R6060 a_3329_8823.n68 a_3329_8823.n67 75.4751
R6061 a_3329_8823.n66 a_3329_8823.n65 75.4751
R6062 a_3329_8823.n15 a_3329_8823.n13 70.8256
R6063 a_3329_8823.n34 a_3329_8823.n32 70.8255
R6064 a_3329_8823.n43 a_3329_8823.n41 70.8255
R6065 a_3329_8823.n24 a_3329_8823.n22 70.8255
R6066 a_3329_8823.n50 a_3329_8823.n49 69.6895
R6067 a_3329_8823.n34 a_3329_8823.n33 69.6895
R6068 a_3329_8823.n36 a_3329_8823.n35 69.6895
R6069 a_3329_8823.n38 a_3329_8823.n37 69.6895
R6070 a_3329_8823.n40 a_3329_8823.n39 69.6895
R6071 a_3329_8823.n43 a_3329_8823.n42 69.6895
R6072 a_3329_8823.n45 a_3329_8823.n44 69.6895
R6073 a_3329_8823.n47 a_3329_8823.n46 69.6895
R6074 a_3329_8823.n31 a_3329_8823.n30 69.6895
R6075 a_3329_8823.n15 a_3329_8823.n14 69.6895
R6076 a_3329_8823.n17 a_3329_8823.n16 69.6895
R6077 a_3329_8823.n19 a_3329_8823.n18 69.6895
R6078 a_3329_8823.n21 a_3329_8823.n20 69.6895
R6079 a_3329_8823.n24 a_3329_8823.n23 69.6895
R6080 a_3329_8823.n26 a_3329_8823.n25 69.6895
R6081 a_3329_8823.n28 a_3329_8823.n27 69.6895
R6082 a_3329_8823.n75 a_3329_8823.t5 17.4005
R6083 a_3329_8823.n75 a_3329_8823.t22 17.4005
R6084 a_3329_8823.n49 a_3329_8823.t73 17.4005
R6085 a_3329_8823.n49 a_3329_8823.t67 17.4005
R6086 a_3329_8823.n32 a_3329_8823.t68 17.4005
R6087 a_3329_8823.n32 a_3329_8823.t77 17.4005
R6088 a_3329_8823.n33 a_3329_8823.t74 17.4005
R6089 a_3329_8823.n33 a_3329_8823.t66 17.4005
R6090 a_3329_8823.n35 a_3329_8823.t46 17.4005
R6091 a_3329_8823.n35 a_3329_8823.t59 17.4005
R6092 a_3329_8823.n37 a_3329_8823.t41 17.4005
R6093 a_3329_8823.n37 a_3329_8823.t42 17.4005
R6094 a_3329_8823.n39 a_3329_8823.t44 17.4005
R6095 a_3329_8823.n39 a_3329_8823.t61 17.4005
R6096 a_3329_8823.n41 a_3329_8823.t49 17.4005
R6097 a_3329_8823.n41 a_3329_8823.t58 17.4005
R6098 a_3329_8823.n42 a_3329_8823.t51 17.4005
R6099 a_3329_8823.n42 a_3329_8823.t79 17.4005
R6100 a_3329_8823.n44 a_3329_8823.t55 17.4005
R6101 a_3329_8823.n44 a_3329_8823.t63 17.4005
R6102 a_3329_8823.n46 a_3329_8823.t54 17.4005
R6103 a_3329_8823.n46 a_3329_8823.t71 17.4005
R6104 a_3329_8823.n30 a_3329_8823.t72 17.4005
R6105 a_3329_8823.n30 a_3329_8823.t60 17.4005
R6106 a_3329_8823.n13 a_3329_8823.t47 17.4005
R6107 a_3329_8823.n13 a_3329_8823.t43 17.4005
R6108 a_3329_8823.n14 a_3329_8823.t64 17.4005
R6109 a_3329_8823.n14 a_3329_8823.t76 17.4005
R6110 a_3329_8823.n16 a_3329_8823.t56 17.4005
R6111 a_3329_8823.n16 a_3329_8823.t65 17.4005
R6112 a_3329_8823.n18 a_3329_8823.t70 17.4005
R6113 a_3329_8823.n18 a_3329_8823.t75 17.4005
R6114 a_3329_8823.n20 a_3329_8823.t40 17.4005
R6115 a_3329_8823.n20 a_3329_8823.t45 17.4005
R6116 a_3329_8823.n22 a_3329_8823.t78 17.4005
R6117 a_3329_8823.n22 a_3329_8823.t50 17.4005
R6118 a_3329_8823.n23 a_3329_8823.t62 17.4005
R6119 a_3329_8823.n23 a_3329_8823.t48 17.4005
R6120 a_3329_8823.n25 a_3329_8823.t69 17.4005
R6121 a_3329_8823.n25 a_3329_8823.t53 17.4005
R6122 a_3329_8823.n27 a_3329_8823.t57 17.4005
R6123 a_3329_8823.n27 a_3329_8823.t52 17.4005
R6124 a_3329_8823.n11 a_3329_8823.t10 17.4005
R6125 a_3329_8823.n11 a_3329_8823.t35 17.4005
R6126 a_3329_8823.n9 a_3329_8823.t21 17.4005
R6127 a_3329_8823.n9 a_3329_8823.t23 17.4005
R6128 a_3329_8823.n7 a_3329_8823.t31 17.4005
R6129 a_3329_8823.n7 a_3329_8823.t16 17.4005
R6130 a_3329_8823.n6 a_3329_8823.t4 17.4005
R6131 a_3329_8823.n6 a_3329_8823.t2 17.4005
R6132 a_3329_8823.n4 a_3329_8823.t34 17.4005
R6133 a_3329_8823.n4 a_3329_8823.t30 17.4005
R6134 a_3329_8823.n3 a_3329_8823.t36 17.4005
R6135 a_3329_8823.n3 a_3329_8823.t27 17.4005
R6136 a_3329_8823.n1 a_3329_8823.t15 17.4005
R6137 a_3329_8823.n1 a_3329_8823.t33 17.4005
R6138 a_3329_8823.n0 a_3329_8823.t24 17.4005
R6139 a_3329_8823.n0 a_3329_8823.t9 17.4005
R6140 a_3329_8823.n56 a_3329_8823.t37 17.4005
R6141 a_3329_8823.n56 a_3329_8823.t20 17.4005
R6142 a_3329_8823.n55 a_3329_8823.t14 17.4005
R6143 a_3329_8823.n55 a_3329_8823.t13 17.4005
R6144 a_3329_8823.n59 a_3329_8823.t26 17.4005
R6145 a_3329_8823.n59 a_3329_8823.t28 17.4005
R6146 a_3329_8823.n58 a_3329_8823.t17 17.4005
R6147 a_3329_8823.n58 a_3329_8823.t7 17.4005
R6148 a_3329_8823.n62 a_3329_8823.t11 17.4005
R6149 a_3329_8823.n62 a_3329_8823.t12 17.4005
R6150 a_3329_8823.n61 a_3329_8823.t3 17.4005
R6151 a_3329_8823.n61 a_3329_8823.t29 17.4005
R6152 a_3329_8823.n69 a_3329_8823.t8 17.4005
R6153 a_3329_8823.n69 a_3329_8823.t1 17.4005
R6154 a_3329_8823.n67 a_3329_8823.t39 17.4005
R6155 a_3329_8823.n67 a_3329_8823.t38 17.4005
R6156 a_3329_8823.n65 a_3329_8823.t18 17.4005
R6157 a_3329_8823.n65 a_3329_8823.t19 17.4005
R6158 a_3329_8823.n64 a_3329_8823.t25 17.4005
R6159 a_3329_8823.n64 a_3329_8823.t6 17.4005
R6160 a_3329_8823.n77 a_3329_8823.t32 17.4005
R6161 a_3329_8823.t0 a_3329_8823.n77 17.4005
R6162 a_3329_8823.n52 a_3329_8823.n51 9.87647
R6163 a_3329_8823.n51 a_3329_8823.n50 2.65128
R6164 a_3329_8823.n48 a_3329_8823.n47 1.78861
R6165 a_3329_8823.n29 a_3329_8823.n28 1.78861
R6166 a_3329_8823.n51 a_3329_8823.n31 1.41089
R6167 a_3329_8823.n40 a_3329_8823.n38 1.14737
R6168 a_3329_8823.n47 a_3329_8823.n45 1.14737
R6169 a_3329_8823.n21 a_3329_8823.n19 1.14737
R6170 a_3329_8823.n28 a_3329_8823.n26 1.14737
R6171 a_3329_8823.n36 a_3329_8823.n34 1.1365
R6172 a_3329_8823.n38 a_3329_8823.n36 1.1365
R6173 a_3329_8823.n45 a_3329_8823.n43 1.1365
R6174 a_3329_8823.n17 a_3329_8823.n15 1.1365
R6175 a_3329_8823.n19 a_3329_8823.n17 1.1365
R6176 a_3329_8823.n26 a_3329_8823.n24 1.1365
R6177 a_3329_8823.n54 a_3329_8823.n2 0.912431
R6178 a_3329_8823.n73 a_3329_8823.n57 0.912431
R6179 a_3329_8823.n71 a_3329_8823.n63 0.912431
R6180 a_3329_8823.n71 a_3329_8823.n70 0.841084
R6181 a_3329_8823.n50 a_3329_8823.n48 0.636437
R6182 a_3329_8823.n31 a_3329_8823.n29 0.636437
R6183 a_3329_8823.n52 a_3329_8823.n12 0.575597
R6184 a_3329_8823.n53 a_3329_8823.n5 0.575597
R6185 a_3329_8823.n72 a_3329_8823.n60 0.575597
R6186 a_3329_8823.n76 a_3329_8823.n74 0.575597
R6187 a_3329_8823.n48 a_3329_8823.n40 0.386435
R6188 a_3329_8823.n29 a_3329_8823.n21 0.386435
R6189 a_3329_8823.n10 a_3329_8823.n8 0.337333
R6190 a_3329_8823.n12 a_3329_8823.n10 0.337333
R6191 a_3329_8823.n68 a_3329_8823.n66 0.337333
R6192 a_3329_8823.n70 a_3329_8823.n68 0.337333
R6193 a_3329_8823.n54 a_3329_8823.n53 0.265986
R6194 a_3329_8823.n74 a_3329_8823.n54 0.265986
R6195 a_3329_8823.n74 a_3329_8823.n73 0.265986
R6196 a_3329_8823.n73 a_3329_8823.n72 0.265986
R6197 a_3329_8823.n72 a_3329_8823.n71 0.265986
R6198 a_3329_8823.n53 a_3329_8823.n52 0.264716
R6199 a_3868_4185.n61 a_3868_4185.n59 70.8256
R6200 a_3868_4185.n2 a_3868_4185.n0 70.8255
R6201 a_3868_4185.n30 a_3868_4185.n28 70.8255
R6202 a_3868_4185.n15 a_3868_4185.n13 70.8255
R6203 a_3868_4185.n46 a_3868_4185.n44 70.8255
R6204 a_3868_4185.n2 a_3868_4185.n1 69.6895
R6205 a_3868_4185.n4 a_3868_4185.n3 69.6895
R6206 a_3868_4185.n6 a_3868_4185.n5 69.6895
R6207 a_3868_4185.n8 a_3868_4185.n7 69.6895
R6208 a_3868_4185.n10 a_3868_4185.n9 69.6895
R6209 a_3868_4185.n12 a_3868_4185.n11 69.6895
R6210 a_3868_4185.n30 a_3868_4185.n29 69.6895
R6211 a_3868_4185.n32 a_3868_4185.n31 69.6895
R6212 a_3868_4185.n34 a_3868_4185.n33 69.6895
R6213 a_3868_4185.n36 a_3868_4185.n35 69.6895
R6214 a_3868_4185.n38 a_3868_4185.n37 69.6895
R6215 a_3868_4185.n40 a_3868_4185.n39 69.6895
R6216 a_3868_4185.n42 a_3868_4185.n41 69.6895
R6217 a_3868_4185.n15 a_3868_4185.n14 69.6895
R6218 a_3868_4185.n17 a_3868_4185.n16 69.6895
R6219 a_3868_4185.n19 a_3868_4185.n18 69.6895
R6220 a_3868_4185.n21 a_3868_4185.n20 69.6895
R6221 a_3868_4185.n23 a_3868_4185.n22 69.6895
R6222 a_3868_4185.n25 a_3868_4185.n24 69.6895
R6223 a_3868_4185.n27 a_3868_4185.n26 69.6895
R6224 a_3868_4185.n46 a_3868_4185.n45 69.6895
R6225 a_3868_4185.n48 a_3868_4185.n47 69.6895
R6226 a_3868_4185.n50 a_3868_4185.n49 69.6895
R6227 a_3868_4185.n52 a_3868_4185.n51 69.6895
R6228 a_3868_4185.n54 a_3868_4185.n53 69.6895
R6229 a_3868_4185.n56 a_3868_4185.n55 69.6895
R6230 a_3868_4185.n58 a_3868_4185.n57 69.6895
R6231 a_3868_4185.n61 a_3868_4185.n60 69.6895
R6232 a_3868_4185.n63 a_3868_4185.n62 69.6895
R6233 a_3868_4185.n65 a_3868_4185.n64 69.6895
R6234 a_3868_4185.n67 a_3868_4185.n66 69.6895
R6235 a_3868_4185.n69 a_3868_4185.n68 69.6895
R6236 a_3868_4185.n71 a_3868_4185.n70 69.6895
R6237 a_3868_4185.n73 a_3868_4185.n72 69.6895
R6238 a_3868_4185.n77 a_3868_4185.n76 69.6895
R6239 a_3868_4185.n0 a_3868_4185.t17 17.4005
R6240 a_3868_4185.n0 a_3868_4185.t16 17.4005
R6241 a_3868_4185.n1 a_3868_4185.t28 17.4005
R6242 a_3868_4185.n1 a_3868_4185.t73 17.4005
R6243 a_3868_4185.n3 a_3868_4185.t62 17.4005
R6244 a_3868_4185.n3 a_3868_4185.t5 17.4005
R6245 a_3868_4185.n5 a_3868_4185.t27 17.4005
R6246 a_3868_4185.n5 a_3868_4185.t70 17.4005
R6247 a_3868_4185.n7 a_3868_4185.t61 17.4005
R6248 a_3868_4185.n7 a_3868_4185.t4 17.4005
R6249 a_3868_4185.n9 a_3868_4185.t11 17.4005
R6250 a_3868_4185.n9 a_3868_4185.t65 17.4005
R6251 a_3868_4185.n11 a_3868_4185.t79 17.4005
R6252 a_3868_4185.n11 a_3868_4185.t31 17.4005
R6253 a_3868_4185.n28 a_3868_4185.t51 17.4005
R6254 a_3868_4185.n28 a_3868_4185.t34 17.4005
R6255 a_3868_4185.n29 a_3868_4185.t55 17.4005
R6256 a_3868_4185.n29 a_3868_4185.t63 17.4005
R6257 a_3868_4185.n31 a_3868_4185.t46 17.4005
R6258 a_3868_4185.n31 a_3868_4185.t25 17.4005
R6259 a_3868_4185.n33 a_3868_4185.t54 17.4005
R6260 a_3868_4185.n33 a_3868_4185.t60 17.4005
R6261 a_3868_4185.n35 a_3868_4185.t45 17.4005
R6262 a_3868_4185.n35 a_3868_4185.t26 17.4005
R6263 a_3868_4185.n37 a_3868_4185.t48 17.4005
R6264 a_3868_4185.n37 a_3868_4185.t76 17.4005
R6265 a_3868_4185.n39 a_3868_4185.t40 17.4005
R6266 a_3868_4185.n39 a_3868_4185.t10 17.4005
R6267 a_3868_4185.n41 a_3868_4185.t44 17.4005
R6268 a_3868_4185.n41 a_3868_4185.t19 17.4005
R6269 a_3868_4185.n13 a_3868_4185.t33 17.4005
R6270 a_3868_4185.n13 a_3868_4185.t1 17.4005
R6271 a_3868_4185.n14 a_3868_4185.t59 17.4005
R6272 a_3868_4185.n14 a_3868_4185.t15 17.4005
R6273 a_3868_4185.n16 a_3868_4185.t22 17.4005
R6274 a_3868_4185.n16 a_3868_4185.t78 17.4005
R6275 a_3868_4185.n18 a_3868_4185.t58 17.4005
R6276 a_3868_4185.n18 a_3868_4185.t14 17.4005
R6277 a_3868_4185.n20 a_3868_4185.t21 17.4005
R6278 a_3868_4185.n20 a_3868_4185.t77 17.4005
R6279 a_3868_4185.n22 a_3868_4185.t74 17.4005
R6280 a_3868_4185.n22 a_3868_4185.t36 17.4005
R6281 a_3868_4185.n24 a_3868_4185.t9 17.4005
R6282 a_3868_4185.n24 a_3868_4185.t67 17.4005
R6283 a_3868_4185.n26 a_3868_4185.t18 17.4005
R6284 a_3868_4185.n26 a_3868_4185.t29 17.4005
R6285 a_3868_4185.n44 a_3868_4185.t13 17.4005
R6286 a_3868_4185.n44 a_3868_4185.t12 17.4005
R6287 a_3868_4185.n45 a_3868_4185.t69 17.4005
R6288 a_3868_4185.n45 a_3868_4185.t24 17.4005
R6289 a_3868_4185.n47 a_3868_4185.t3 17.4005
R6290 a_3868_4185.n47 a_3868_4185.t57 17.4005
R6291 a_3868_4185.n49 a_3868_4185.t68 17.4005
R6292 a_3868_4185.n49 a_3868_4185.t23 17.4005
R6293 a_3868_4185.n51 a_3868_4185.t2 17.4005
R6294 a_3868_4185.n51 a_3868_4185.t56 17.4005
R6295 a_3868_4185.n53 a_3868_4185.t64 17.4005
R6296 a_3868_4185.n53 a_3868_4185.t8 17.4005
R6297 a_3868_4185.n55 a_3868_4185.t30 17.4005
R6298 a_3868_4185.n55 a_3868_4185.t75 17.4005
R6299 a_3868_4185.n57 a_3868_4185.t38 17.4005
R6300 a_3868_4185.n57 a_3868_4185.t37 17.4005
R6301 a_3868_4185.n59 a_3868_4185.t35 17.4005
R6302 a_3868_4185.n59 a_3868_4185.t53 17.4005
R6303 a_3868_4185.n60 a_3868_4185.t7 17.4005
R6304 a_3868_4185.n60 a_3868_4185.t42 17.4005
R6305 a_3868_4185.n62 a_3868_4185.t72 17.4005
R6306 a_3868_4185.n62 a_3868_4185.t50 17.4005
R6307 a_3868_4185.n64 a_3868_4185.t6 17.4005
R6308 a_3868_4185.n64 a_3868_4185.t41 17.4005
R6309 a_3868_4185.n66 a_3868_4185.t71 17.4005
R6310 a_3868_4185.n66 a_3868_4185.t49 17.4005
R6311 a_3868_4185.n68 a_3868_4185.t32 17.4005
R6312 a_3868_4185.n68 a_3868_4185.t52 17.4005
R6313 a_3868_4185.n70 a_3868_4185.t66 17.4005
R6314 a_3868_4185.n70 a_3868_4185.t43 17.4005
R6315 a_3868_4185.n72 a_3868_4185.t20 17.4005
R6316 a_3868_4185.n72 a_3868_4185.t47 17.4005
R6317 a_3868_4185.n77 a_3868_4185.t0 17.4005
R6318 a_3868_4185.t39 a_3868_4185.n77 17.4005
R6319 a_3868_4185.n43 a_3868_4185.n42 2.29404
R6320 a_3868_4185.n74 a_3868_4185.n73 2.29404
R6321 a_3868_4185.n75 a_3868_4185.n43 1.40267
R6322 a_3868_4185.n75 a_3868_4185.n74 1.40267
R6323 a_3868_4185.n32 a_3868_4185.n30 1.1365
R6324 a_3868_4185.n34 a_3868_4185.n32 1.1365
R6325 a_3868_4185.n36 a_3868_4185.n34 1.1365
R6326 a_3868_4185.n38 a_3868_4185.n36 1.1365
R6327 a_3868_4185.n40 a_3868_4185.n38 1.1365
R6328 a_3868_4185.n42 a_3868_4185.n40 1.1365
R6329 a_3868_4185.n17 a_3868_4185.n15 1.1365
R6330 a_3868_4185.n19 a_3868_4185.n17 1.1365
R6331 a_3868_4185.n21 a_3868_4185.n19 1.1365
R6332 a_3868_4185.n23 a_3868_4185.n21 1.1365
R6333 a_3868_4185.n25 a_3868_4185.n23 1.1365
R6334 a_3868_4185.n27 a_3868_4185.n25 1.1365
R6335 a_3868_4185.n48 a_3868_4185.n46 1.1365
R6336 a_3868_4185.n50 a_3868_4185.n48 1.1365
R6337 a_3868_4185.n52 a_3868_4185.n50 1.1365
R6338 a_3868_4185.n54 a_3868_4185.n52 1.1365
R6339 a_3868_4185.n56 a_3868_4185.n54 1.1365
R6340 a_3868_4185.n58 a_3868_4185.n56 1.1365
R6341 a_3868_4185.n63 a_3868_4185.n61 1.1365
R6342 a_3868_4185.n65 a_3868_4185.n63 1.1365
R6343 a_3868_4185.n67 a_3868_4185.n65 1.1365
R6344 a_3868_4185.n69 a_3868_4185.n67 1.1365
R6345 a_3868_4185.n71 a_3868_4185.n69 1.1365
R6346 a_3868_4185.n73 a_3868_4185.n71 1.1365
R6347 a_3868_4185.n4 a_3868_4185.n2 1.1365
R6348 a_3868_4185.n6 a_3868_4185.n4 1.1365
R6349 a_3868_4185.n8 a_3868_4185.n6 1.1365
R6350 a_3868_4185.n10 a_3868_4185.n8 1.1365
R6351 a_3868_4185.n12 a_3868_4185.n10 1.1365
R6352 a_3868_4185.n76 a_3868_4185.n12 1.1365
R6353 a_3868_4185.n43 a_3868_4185.n27 0.89187
R6354 a_3868_4185.n74 a_3868_4185.n58 0.89187
R6355 a_3868_4185.n76 a_3868_4185.n75 0.89187
R6356 VOUT.n15 VOUT.n13 204.214
R6357 VOUT.n2 VOUT.n0 204.214
R6358 VOUT.n2 VOUT.n1 203.03
R6359 VOUT.n4 VOUT.n3 203.03
R6360 VOUT.n6 VOUT.n5 203.03
R6361 VOUT.n8 VOUT.n7 203.03
R6362 VOUT.n10 VOUT.n9 203.03
R6363 VOUT.n12 VOUT.n11 203.03
R6364 VOUT.n15 VOUT.n14 203.03
R6365 VOUT.n17 VOUT.n16 203.03
R6366 VOUT.n19 VOUT.n18 203.03
R6367 VOUT.n21 VOUT.n20 203.03
R6368 VOUT.n23 VOUT.n22 203.03
R6369 VOUT.n25 VOUT.n24 203.03
R6370 VOUT.n68 VOUT.n66 76.1487
R6371 VOUT.n63 VOUT.n61 76.1487
R6372 VOUT.n58 VOUT.n56 76.1487
R6373 VOUT.n53 VOUT.n51 76.1487
R6374 VOUT.n48 VOUT.n46 76.1487
R6375 VOUT.n43 VOUT.n41 76.1487
R6376 VOUT.n38 VOUT.n36 76.1487
R6377 VOUT.n33 VOUT.n31 76.1487
R6378 VOUT.n73 VOUT.n71 75.8119
R6379 VOUT.n28 VOUT.n26 75.8119
R6380 VOUT.n75 VOUT.n74 75.4751
R6381 VOUT.n73 VOUT.n72 75.4751
R6382 VOUT.n70 VOUT.n69 75.4751
R6383 VOUT.n68 VOUT.n67 75.4751
R6384 VOUT.n65 VOUT.n64 75.4751
R6385 VOUT.n63 VOUT.n62 75.4751
R6386 VOUT.n60 VOUT.n59 75.4751
R6387 VOUT.n58 VOUT.n57 75.4751
R6388 VOUT.n55 VOUT.n54 75.4751
R6389 VOUT.n53 VOUT.n52 75.4751
R6390 VOUT.n50 VOUT.n49 75.4751
R6391 VOUT.n48 VOUT.n47 75.4751
R6392 VOUT.n45 VOUT.n44 75.4751
R6393 VOUT.n43 VOUT.n42 75.4751
R6394 VOUT.n40 VOUT.n39 75.4751
R6395 VOUT.n38 VOUT.n37 75.4751
R6396 VOUT.n35 VOUT.n34 75.4751
R6397 VOUT.n33 VOUT.n32 75.4751
R6398 VOUT.n30 VOUT.n29 75.4751
R6399 VOUT.n28 VOUT.n27 75.4751
R6400 VOUT.n0 VOUT.t65 28.5655
R6401 VOUT.n0 VOUT.t69 28.5655
R6402 VOUT.n1 VOUT.t75 28.5655
R6403 VOUT.n1 VOUT.t73 28.5655
R6404 VOUT.n3 VOUT.t64 28.5655
R6405 VOUT.n3 VOUT.t63 28.5655
R6406 VOUT.n5 VOUT.t83 28.5655
R6407 VOUT.n5 VOUT.t80 28.5655
R6408 VOUT.n7 VOUT.t86 28.5655
R6409 VOUT.n7 VOUT.t79 28.5655
R6410 VOUT.n9 VOUT.t67 28.5655
R6411 VOUT.n9 VOUT.t81 28.5655
R6412 VOUT.n11 VOUT.t71 28.5655
R6413 VOUT.n11 VOUT.t85 28.5655
R6414 VOUT.n13 VOUT.t76 28.5655
R6415 VOUT.n13 VOUT.t74 28.5655
R6416 VOUT.n14 VOUT.t70 28.5655
R6417 VOUT.n14 VOUT.t82 28.5655
R6418 VOUT.n16 VOUT.t87 28.5655
R6419 VOUT.n16 VOUT.t66 28.5655
R6420 VOUT.n18 VOUT.t62 28.5655
R6421 VOUT.n18 VOUT.t60 28.5655
R6422 VOUT.n20 VOUT.t61 28.5655
R6423 VOUT.n20 VOUT.t88 28.5655
R6424 VOUT.n22 VOUT.t84 28.5655
R6425 VOUT.n22 VOUT.t68 28.5655
R6426 VOUT.n24 VOUT.t77 28.5655
R6427 VOUT.n24 VOUT.t72 28.5655
R6428 VOUT.n86 VOUT.n85 17.5151
R6429 VOUT.n74 VOUT.t45 17.4005
R6430 VOUT.n74 VOUT.t25 17.4005
R6431 VOUT.n72 VOUT.t48 17.4005
R6432 VOUT.n72 VOUT.t46 17.4005
R6433 VOUT.n71 VOUT.t13 17.4005
R6434 VOUT.n71 VOUT.t56 17.4005
R6435 VOUT.n69 VOUT.t18 17.4005
R6436 VOUT.n69 VOUT.t41 17.4005
R6437 VOUT.n67 VOUT.t55 17.4005
R6438 VOUT.n67 VOUT.t51 17.4005
R6439 VOUT.n66 VOUT.t42 17.4005
R6440 VOUT.n66 VOUT.t35 17.4005
R6441 VOUT.n64 VOUT.t52 17.4005
R6442 VOUT.n64 VOUT.t54 17.4005
R6443 VOUT.n62 VOUT.t2 17.4005
R6444 VOUT.n62 VOUT.t26 17.4005
R6445 VOUT.n61 VOUT.t39 17.4005
R6446 VOUT.n61 VOUT.t34 17.4005
R6447 VOUT.n59 VOUT.t47 17.4005
R6448 VOUT.n59 VOUT.t38 17.4005
R6449 VOUT.n57 VOUT.t43 17.4005
R6450 VOUT.n57 VOUT.t44 17.4005
R6451 VOUT.n56 VOUT.t58 17.4005
R6452 VOUT.n56 VOUT.t16 17.4005
R6453 VOUT.n54 VOUT.t15 17.4005
R6454 VOUT.n54 VOUT.t40 17.4005
R6455 VOUT.n52 VOUT.t22 17.4005
R6456 VOUT.n52 VOUT.t10 17.4005
R6457 VOUT.n51 VOUT.t31 17.4005
R6458 VOUT.n51 VOUT.t33 17.4005
R6459 VOUT.n49 VOUT.t9 17.4005
R6460 VOUT.n49 VOUT.t14 17.4005
R6461 VOUT.n47 VOUT.t21 17.4005
R6462 VOUT.n47 VOUT.t0 17.4005
R6463 VOUT.n46 VOUT.t20 17.4005
R6464 VOUT.n46 VOUT.t8 17.4005
R6465 VOUT.n44 VOUT.t12 17.4005
R6466 VOUT.n44 VOUT.t36 17.4005
R6467 VOUT.n42 VOUT.t32 17.4005
R6468 VOUT.n42 VOUT.t1 17.4005
R6469 VOUT.n41 VOUT.t27 17.4005
R6470 VOUT.n41 VOUT.t49 17.4005
R6471 VOUT.n39 VOUT.t3 17.4005
R6472 VOUT.n39 VOUT.t17 17.4005
R6473 VOUT.n37 VOUT.t53 17.4005
R6474 VOUT.n37 VOUT.t6 17.4005
R6475 VOUT.n36 VOUT.t11 17.4005
R6476 VOUT.n36 VOUT.t19 17.4005
R6477 VOUT.n34 VOUT.t5 17.4005
R6478 VOUT.n34 VOUT.t37 17.4005
R6479 VOUT.n32 VOUT.t4 17.4005
R6480 VOUT.n32 VOUT.t7 17.4005
R6481 VOUT.n31 VOUT.t59 17.4005
R6482 VOUT.n31 VOUT.t28 17.4005
R6483 VOUT.n29 VOUT.t29 17.4005
R6484 VOUT.n29 VOUT.t24 17.4005
R6485 VOUT.n27 VOUT.t50 17.4005
R6486 VOUT.n27 VOUT.t30 17.4005
R6487 VOUT.n26 VOUT.t57 17.4005
R6488 VOUT.n26 VOUT.t23 17.4005
R6489 VOUT.n85 VOUT.n84 16.8905
R6490 VOUT VOUT.n87 13.3103
R6491 VOUT.n76 VOUT.n75 1.51348
R6492 VOUT.n87 VOUT.n86 1.40267
R6493 VOUT.n87 VOUT.n12 1.40003
R6494 VOUT.n86 VOUT.n25 1.40003
R6495 VOUT.n4 VOUT.n2 1.18544
R6496 VOUT.n6 VOUT.n4 1.18544
R6497 VOUT.n8 VOUT.n6 1.18544
R6498 VOUT.n10 VOUT.n8 1.18544
R6499 VOUT.n12 VOUT.n10 1.18544
R6500 VOUT.n17 VOUT.n15 1.18544
R6501 VOUT.n19 VOUT.n17 1.18544
R6502 VOUT.n21 VOUT.n19 1.18544
R6503 VOUT.n23 VOUT.n21 1.18544
R6504 VOUT.n25 VOUT.n23 1.18544
R6505 VOUT.n76 VOUT.n70 0.912431
R6506 VOUT.n78 VOUT.n60 0.912431
R6507 VOUT.n80 VOUT.n50 0.912431
R6508 VOUT.n82 VOUT.n40 0.912431
R6509 VOUT.n84 VOUT.n30 0.912431
R6510 VOUT.n70 VOUT.n68 0.674167
R6511 VOUT.n65 VOUT.n63 0.674167
R6512 VOUT.n60 VOUT.n58 0.674167
R6513 VOUT.n55 VOUT.n53 0.674167
R6514 VOUT.n50 VOUT.n48 0.674167
R6515 VOUT.n45 VOUT.n43 0.674167
R6516 VOUT.n40 VOUT.n38 0.674167
R6517 VOUT.n35 VOUT.n33 0.674167
R6518 VOUT.n77 VOUT.n65 0.575597
R6519 VOUT.n79 VOUT.n55 0.575597
R6520 VOUT.n81 VOUT.n45 0.575597
R6521 VOUT.n83 VOUT.n35 0.575597
R6522 VOUT.n75 VOUT.n73 0.337333
R6523 VOUT.n30 VOUT.n28 0.337333
R6524 VOUT.n77 VOUT.n76 0.265986
R6525 VOUT.n78 VOUT.n77 0.265986
R6526 VOUT.n79 VOUT.n78 0.265986
R6527 VOUT.n80 VOUT.n79 0.265986
R6528 VOUT.n81 VOUT.n80 0.265986
R6529 VOUT.n82 VOUT.n81 0.265986
R6530 VOUT.n83 VOUT.n82 0.265986
R6531 VOUT.n84 VOUT.n83 0.265986
R6532 VOUT.n85 VOUT.t78 0.0115332
R6533 a_n1962_4406.n21 a_n1962_4406.n19 70.8256
R6534 a_n1962_4406.n115 a_n1962_4406.n113 70.8255
R6535 a_n1962_4406.n2 a_n1962_4406.n0 70.8255
R6536 a_n1962_4406.n8 a_n1962_4406.n6 70.8255
R6537 a_n1962_4406.n58 a_n1962_4406.n56 70.8255
R6538 a_n1962_4406.n25 a_n1962_4406.n23 70.8255
R6539 a_n1962_4406.n39 a_n1962_4406.n37 70.8255
R6540 a_n1962_4406.n5 a_n1962_4406.n3 70.8255
R6541 a_n1962_4406.n98 a_n1962_4406.n96 70.8255
R6542 a_n1962_4406.n79 a_n1962_4406.n77 70.8255
R6543 a_n1962_4406.n83 a_n1962_4406.n81 70.8255
R6544 a_n1962_4406.n48 a_n1962_4406.n36 70.2276
R6545 a_n1962_4406.n52 a_n1962_4406.n22 70.1244
R6546 a_n1962_4406.n92 a_n1962_4406.n80 70.1054
R6547 a_n1962_4406.n110 a_n1962_4406.n109 69.6895
R6548 a_n1962_4406.n112 a_n1962_4406.n111 69.6895
R6549 a_n1962_4406.n119 a_n1962_4406.n118 69.6895
R6550 a_n1962_4406.n117 a_n1962_4406.n116 69.6895
R6551 a_n1962_4406.n115 a_n1962_4406.n114 69.6895
R6552 a_n1962_4406.n76 a_n1962_4406.n75 69.6895
R6553 a_n1962_4406.n2 a_n1962_4406.n1 69.6895
R6554 a_n1962_4406.n72 a_n1962_4406.n71 69.6895
R6555 a_n1962_4406.n18 a_n1962_4406.n17 69.6895
R6556 a_n1962_4406.n16 a_n1962_4406.n15 69.6895
R6557 a_n1962_4406.n14 a_n1962_4406.n13 69.6895
R6558 a_n1962_4406.n12 a_n1962_4406.n11 69.6895
R6559 a_n1962_4406.n10 a_n1962_4406.n9 69.6895
R6560 a_n1962_4406.n8 a_n1962_4406.n7 69.6895
R6561 a_n1962_4406.n68 a_n1962_4406.n67 69.6895
R6562 a_n1962_4406.n66 a_n1962_4406.n65 69.6895
R6563 a_n1962_4406.n64 a_n1962_4406.n63 69.6895
R6564 a_n1962_4406.n62 a_n1962_4406.n61 69.6895
R6565 a_n1962_4406.n60 a_n1962_4406.n59 69.6895
R6566 a_n1962_4406.n58 a_n1962_4406.n57 69.6895
R6567 a_n1962_4406.n55 a_n1962_4406.n54 69.6895
R6568 a_n1962_4406.n21 a_n1962_4406.n20 69.6895
R6569 a_n1962_4406.n51 a_n1962_4406.n50 69.6895
R6570 a_n1962_4406.n35 a_n1962_4406.n34 69.6895
R6571 a_n1962_4406.n33 a_n1962_4406.n32 69.6895
R6572 a_n1962_4406.n31 a_n1962_4406.n30 69.6895
R6573 a_n1962_4406.n29 a_n1962_4406.n28 69.6895
R6574 a_n1962_4406.n27 a_n1962_4406.n26 69.6895
R6575 a_n1962_4406.n25 a_n1962_4406.n24 69.6895
R6576 a_n1962_4406.n47 a_n1962_4406.n46 69.6895
R6577 a_n1962_4406.n45 a_n1962_4406.n44 69.6895
R6578 a_n1962_4406.n43 a_n1962_4406.n42 69.6895
R6579 a_n1962_4406.n41 a_n1962_4406.n40 69.6895
R6580 a_n1962_4406.n39 a_n1962_4406.n38 69.6895
R6581 a_n1962_4406.n5 a_n1962_4406.n4 69.6895
R6582 a_n1962_4406.n106 a_n1962_4406.n105 69.6895
R6583 a_n1962_4406.n104 a_n1962_4406.n103 69.6895
R6584 a_n1962_4406.n102 a_n1962_4406.n101 69.6895
R6585 a_n1962_4406.n100 a_n1962_4406.n99 69.6895
R6586 a_n1962_4406.n98 a_n1962_4406.n97 69.6895
R6587 a_n1962_4406.n95 a_n1962_4406.n94 69.6895
R6588 a_n1962_4406.n79 a_n1962_4406.n78 69.6895
R6589 a_n1962_4406.n91 a_n1962_4406.n90 69.6895
R6590 a_n1962_4406.n89 a_n1962_4406.n88 69.6895
R6591 a_n1962_4406.n87 a_n1962_4406.n86 69.6895
R6592 a_n1962_4406.n85 a_n1962_4406.n84 69.6895
R6593 a_n1962_4406.n83 a_n1962_4406.n82 69.6895
R6594 a_n1962_4406.n121 a_n1962_4406.n120 69.6895
R6595 a_n1962_4406.n109 a_n1962_4406.t102 17.4005
R6596 a_n1962_4406.n109 a_n1962_4406.t13 17.4005
R6597 a_n1962_4406.n111 a_n1962_4406.t2 17.4005
R6598 a_n1962_4406.n111 a_n1962_4406.t112 17.4005
R6599 a_n1962_4406.n118 a_n1962_4406.t47 17.4005
R6600 a_n1962_4406.n118 a_n1962_4406.t99 17.4005
R6601 a_n1962_4406.n116 a_n1962_4406.t88 17.4005
R6602 a_n1962_4406.n116 a_n1962_4406.t58 17.4005
R6603 a_n1962_4406.n114 a_n1962_4406.t46 17.4005
R6604 a_n1962_4406.n114 a_n1962_4406.t98 17.4005
R6605 a_n1962_4406.n113 a_n1962_4406.t60 17.4005
R6606 a_n1962_4406.n113 a_n1962_4406.t45 17.4005
R6607 a_n1962_4406.n75 a_n1962_4406.t20 17.4005
R6608 a_n1962_4406.n75 a_n1962_4406.t80 17.4005
R6609 a_n1962_4406.n0 a_n1962_4406.t22 17.4005
R6610 a_n1962_4406.n0 a_n1962_4406.t3 17.4005
R6611 a_n1962_4406.n1 a_n1962_4406.t115 17.4005
R6612 a_n1962_4406.n1 a_n1962_4406.t30 17.4005
R6613 a_n1962_4406.n71 a_n1962_4406.t119 17.4005
R6614 a_n1962_4406.n71 a_n1962_4406.t56 17.4005
R6615 a_n1962_4406.n17 a_n1962_4406.t10 17.4005
R6616 a_n1962_4406.n17 a_n1962_4406.t86 17.4005
R6617 a_n1962_4406.n15 a_n1962_4406.t103 17.4005
R6618 a_n1962_4406.n15 a_n1962_4406.t37 17.4005
R6619 a_n1962_4406.n13 a_n1962_4406.t49 17.4005
R6620 a_n1962_4406.n13 a_n1962_4406.t117 17.4005
R6621 a_n1962_4406.n11 a_n1962_4406.t91 17.4005
R6622 a_n1962_4406.n11 a_n1962_4406.t16 17.4005
R6623 a_n1962_4406.n9 a_n1962_4406.t48 17.4005
R6624 a_n1962_4406.n9 a_n1962_4406.t116 17.4005
R6625 a_n1962_4406.n7 a_n1962_4406.t90 17.4005
R6626 a_n1962_4406.n7 a_n1962_4406.t15 17.4005
R6627 a_n1962_4406.n6 a_n1962_4406.t31 17.4005
R6628 a_n1962_4406.n6 a_n1962_4406.t33 17.4005
R6629 a_n1962_4406.n67 a_n1962_4406.t121 17.4005
R6630 a_n1962_4406.n67 a_n1962_4406.t11 17.4005
R6631 a_n1962_4406.n65 a_n1962_4406.t26 17.4005
R6632 a_n1962_4406.n65 a_n1962_4406.t106 17.4005
R6633 a_n1962_4406.n63 a_n1962_4406.t105 17.4005
R6634 a_n1962_4406.n63 a_n1962_4406.t51 17.4005
R6635 a_n1962_4406.n61 a_n1962_4406.t5 17.4005
R6636 a_n1962_4406.n61 a_n1962_4406.t93 17.4005
R6637 a_n1962_4406.n59 a_n1962_4406.t104 17.4005
R6638 a_n1962_4406.n59 a_n1962_4406.t50 17.4005
R6639 a_n1962_4406.n57 a_n1962_4406.t4 17.4005
R6640 a_n1962_4406.n57 a_n1962_4406.t92 17.4005
R6641 a_n1962_4406.n56 a_n1962_4406.t24 17.4005
R6642 a_n1962_4406.n56 a_n1962_4406.t32 17.4005
R6643 a_n1962_4406.n54 a_n1962_4406.t41 17.4005
R6644 a_n1962_4406.n54 a_n1962_4406.t120 17.4005
R6645 a_n1962_4406.n19 a_n1962_4406.t42 17.4005
R6646 a_n1962_4406.n19 a_n1962_4406.t79 17.4005
R6647 a_n1962_4406.n20 a_n1962_4406.t87 17.4005
R6648 a_n1962_4406.n20 a_n1962_4406.t27 17.4005
R6649 a_n1962_4406.n50 a_n1962_4406.t111 17.4005
R6650 a_n1962_4406.n50 a_n1962_4406.t43 17.4005
R6651 a_n1962_4406.n34 a_n1962_4406.t55 17.4005
R6652 a_n1962_4406.n34 a_n1962_4406.t122 17.4005
R6653 a_n1962_4406.n32 a_n1962_4406.t94 17.4005
R6654 a_n1962_4406.n32 a_n1962_4406.t28 17.4005
R6655 a_n1962_4406.n30 a_n1962_4406.t35 17.4005
R6656 a_n1962_4406.n30 a_n1962_4406.t108 17.4005
R6657 a_n1962_4406.n28 a_n1962_4406.t82 17.4005
R6658 a_n1962_4406.n28 a_n1962_4406.t7 17.4005
R6659 a_n1962_4406.n26 a_n1962_4406.t34 17.4005
R6660 a_n1962_4406.n26 a_n1962_4406.t107 17.4005
R6661 a_n1962_4406.n24 a_n1962_4406.t81 17.4005
R6662 a_n1962_4406.n24 a_n1962_4406.t6 17.4005
R6663 a_n1962_4406.n23 a_n1962_4406.t23 17.4005
R6664 a_n1962_4406.n23 a_n1962_4406.t68 17.4005
R6665 a_n1962_4406.n46 a_n1962_4406.t123 17.4005
R6666 a_n1962_4406.n46 a_n1962_4406.t69 17.4005
R6667 a_n1962_4406.n44 a_n1962_4406.t29 17.4005
R6668 a_n1962_4406.n44 a_n1962_4406.t77 17.4005
R6669 a_n1962_4406.n42 a_n1962_4406.t110 17.4005
R6670 a_n1962_4406.n42 a_n1962_4406.t62 17.4005
R6671 a_n1962_4406.n40 a_n1962_4406.t9 17.4005
R6672 a_n1962_4406.n40 a_n1962_4406.t73 17.4005
R6673 a_n1962_4406.n38 a_n1962_4406.t109 17.4005
R6674 a_n1962_4406.n38 a_n1962_4406.t61 17.4005
R6675 a_n1962_4406.n37 a_n1962_4406.t8 17.4005
R6676 a_n1962_4406.n37 a_n1962_4406.t72 17.4005
R6677 a_n1962_4406.n36 a_n1962_4406.t44 17.4005
R6678 a_n1962_4406.n36 a_n1962_4406.t65 17.4005
R6679 a_n1962_4406.n22 a_n1962_4406.t12 17.4005
R6680 a_n1962_4406.n22 a_n1962_4406.t66 17.4005
R6681 a_n1962_4406.n3 a_n1962_4406.t54 17.4005
R6682 a_n1962_4406.n3 a_n1962_4406.t57 17.4005
R6683 a_n1962_4406.n4 a_n1962_4406.t25 17.4005
R6684 a_n1962_4406.n4 a_n1962_4406.t96 17.4005
R6685 a_n1962_4406.n105 a_n1962_4406.t38 17.4005
R6686 a_n1962_4406.n105 a_n1962_4406.t118 17.4005
R6687 a_n1962_4406.n103 a_n1962_4406.t83 17.4005
R6688 a_n1962_4406.n103 a_n1962_4406.t18 17.4005
R6689 a_n1962_4406.n101 a_n1962_4406.t17 17.4005
R6690 a_n1962_4406.n101 a_n1962_4406.t101 17.4005
R6691 a_n1962_4406.n99 a_n1962_4406.t113 17.4005
R6692 a_n1962_4406.n99 a_n1962_4406.t1 17.4005
R6693 a_n1962_4406.n97 a_n1962_4406.t14 17.4005
R6694 a_n1962_4406.n97 a_n1962_4406.t100 17.4005
R6695 a_n1962_4406.n96 a_n1962_4406.t76 17.4005
R6696 a_n1962_4406.n96 a_n1962_4406.t0 17.4005
R6697 a_n1962_4406.n94 a_n1962_4406.t95 17.4005
R6698 a_n1962_4406.n94 a_n1962_4406.t36 17.4005
R6699 a_n1962_4406.n77 a_n1962_4406.t70 17.4005
R6700 a_n1962_4406.n77 a_n1962_4406.t39 17.4005
R6701 a_n1962_4406.n78 a_n1962_4406.t52 17.4005
R6702 a_n1962_4406.n78 a_n1962_4406.t84 17.4005
R6703 a_n1962_4406.n90 a_n1962_4406.t67 17.4005
R6704 a_n1962_4406.n90 a_n1962_4406.t97 17.4005
R6705 a_n1962_4406.n88 a_n1962_4406.t71 17.4005
R6706 a_n1962_4406.n88 a_n1962_4406.t40 17.4005
R6707 a_n1962_4406.n86 a_n1962_4406.t78 17.4005
R6708 a_n1962_4406.n86 a_n1962_4406.t85 17.4005
R6709 a_n1962_4406.n84 a_n1962_4406.t64 17.4005
R6710 a_n1962_4406.n84 a_n1962_4406.t21 17.4005
R6711 a_n1962_4406.n82 a_n1962_4406.t74 17.4005
R6712 a_n1962_4406.n82 a_n1962_4406.t114 17.4005
R6713 a_n1962_4406.n81 a_n1962_4406.t63 17.4005
R6714 a_n1962_4406.n81 a_n1962_4406.t19 17.4005
R6715 a_n1962_4406.n80 a_n1962_4406.t75 17.4005
R6716 a_n1962_4406.n80 a_n1962_4406.t53 17.4005
R6717 a_n1962_4406.n121 a_n1962_4406.t89 17.4005
R6718 a_n1962_4406.t59 a_n1962_4406.n121 17.4005
R6719 a_n1962_4406.n49 a_n1962_4406.n48 1.40267
R6720 a_n1962_4406.n53 a_n1962_4406.n52 1.40267
R6721 a_n1962_4406.n70 a_n1962_4406.n69 1.40267
R6722 a_n1962_4406.n74 a_n1962_4406.n73 1.40267
R6723 a_n1962_4406.n93 a_n1962_4406.n92 1.40267
R6724 a_n1962_4406.n108 a_n1962_4406.n107 1.40267
R6725 a_n1962_4406.n18 a_n1962_4406.n16 1.1365
R6726 a_n1962_4406.n16 a_n1962_4406.n14 1.1365
R6727 a_n1962_4406.n14 a_n1962_4406.n12 1.1365
R6728 a_n1962_4406.n12 a_n1962_4406.n10 1.1365
R6729 a_n1962_4406.n10 a_n1962_4406.n8 1.1365
R6730 a_n1962_4406.n35 a_n1962_4406.n33 1.1365
R6731 a_n1962_4406.n33 a_n1962_4406.n31 1.1365
R6732 a_n1962_4406.n31 a_n1962_4406.n29 1.1365
R6733 a_n1962_4406.n29 a_n1962_4406.n27 1.1365
R6734 a_n1962_4406.n27 a_n1962_4406.n25 1.1365
R6735 a_n1962_4406.n47 a_n1962_4406.n45 1.1365
R6736 a_n1962_4406.n45 a_n1962_4406.n43 1.1365
R6737 a_n1962_4406.n43 a_n1962_4406.n41 1.1365
R6738 a_n1962_4406.n41 a_n1962_4406.n39 1.1365
R6739 a_n1962_4406.n68 a_n1962_4406.n66 1.1365
R6740 a_n1962_4406.n66 a_n1962_4406.n64 1.1365
R6741 a_n1962_4406.n64 a_n1962_4406.n62 1.1365
R6742 a_n1962_4406.n62 a_n1962_4406.n60 1.1365
R6743 a_n1962_4406.n60 a_n1962_4406.n58 1.1365
R6744 a_n1962_4406.n91 a_n1962_4406.n89 1.1365
R6745 a_n1962_4406.n89 a_n1962_4406.n87 1.1365
R6746 a_n1962_4406.n87 a_n1962_4406.n85 1.1365
R6747 a_n1962_4406.n85 a_n1962_4406.n83 1.1365
R6748 a_n1962_4406.n106 a_n1962_4406.n104 1.1365
R6749 a_n1962_4406.n104 a_n1962_4406.n102 1.1365
R6750 a_n1962_4406.n102 a_n1962_4406.n100 1.1365
R6751 a_n1962_4406.n100 a_n1962_4406.n98 1.1365
R6752 a_n1962_4406.n112 a_n1962_4406.n110 1.1365
R6753 a_n1962_4406.n120 a_n1962_4406.n112 1.1365
R6754 a_n1962_4406.n120 a_n1962_4406.n119 1.1365
R6755 a_n1962_4406.n119 a_n1962_4406.n117 1.1365
R6756 a_n1962_4406.n117 a_n1962_4406.n115 1.1365
R6757 a_n1962_4406.n92 a_n1962_4406.n91 0.595676
R6758 a_n1962_4406.n95 a_n1962_4406.n93 0.595676
R6759 a_n1962_4406.n73 a_n1962_4406.n72 0.582089
R6760 a_n1962_4406.n76 a_n1962_4406.n74 0.582089
R6761 a_n1962_4406.n108 a_n1962_4406.n76 0.582087
R6762 a_n1962_4406.n107 a_n1962_4406.n95 0.582087
R6763 a_n1962_4406.n52 a_n1962_4406.n51 0.576654
R6764 a_n1962_4406.n55 a_n1962_4406.n53 0.576654
R6765 a_n1962_4406.n69 a_n1962_4406.n55 0.5685
R6766 a_n1962_4406.n72 a_n1962_4406.n70 0.5685
R6767 a_n1962_4406.n51 a_n1962_4406.n49 0.538609
R6768 a_n1962_4406.n49 a_n1962_4406.n35 0.473394
R6769 a_n1962_4406.n48 a_n1962_4406.n47 0.473394
R6770 a_n1962_4406.n70 a_n1962_4406.n18 0.443502
R6771 a_n1962_4406.n69 a_n1962_4406.n68 0.443502
R6772 a_n1962_4406.n53 a_n1962_4406.n21 0.435348
R6773 a_n1962_4406.n107 a_n1962_4406.n106 0.429915
R6774 a_n1962_4406.n110 a_n1962_4406.n108 0.429915
R6775 a_n1962_4406.n74 a_n1962_4406.n2 0.429914
R6776 a_n1962_4406.n73 a_n1962_4406.n5 0.429914
R6777 a_n1962_4406.n93 a_n1962_4406.n79 0.416327
R6778 VP.n0 VP.t14 118.507
R6779 VP.n1 VP.t12 117.266
R6780 VP.n3 VP.t11 117.266
R6781 VP.n7 VP.t0 117.266
R6782 VP.n9 VP.t9 117.266
R6783 VP.n13 VP.t5 117.266
R6784 VP.n0 VP.t2 116.647
R6785 VP.n1 VP.t4 116.647
R6786 VP.n3 VP.t8 116.647
R6787 VP.n4 VP.t13 116.647
R6788 VP.n5 VP.t1 116.647
R6789 VP.n7 VP.t10 116.647
R6790 VP.n9 VP.t15 116.647
R6791 VP.n10 VP.t7 116.647
R6792 VP.n11 VP.t6 116.647
R6793 VP.n13 VP.t3 116.647
R6794 VP VP.n14 29.6934
R6795 VP.n2 VP.n0 3.71637
R6796 VP.n2 VP.n1 3.32392
R6797 VP.n8 VP.n7 3.32392
R6798 VP.n14 VP.n13 3.32392
R6799 VP.n6 VP.n5 2.08353
R6800 VP.n12 VP.n11 2.08353
R6801 VP.n4 VP.n3 1.85887
R6802 VP.n10 VP.n9 1.85887
R6803 VP.n6 VP.n2 1.00593
R6804 VP.n8 VP.n6 0.995065
R6805 VP.n12 VP.n8 0.995065
R6806 VP.n14 VP.n12 0.995065
R6807 VP.n5 VP.n4 0.618487
R6808 VP.n11 VP.n10 0.618487
R6809 a_n735_8972.n50 a_n735_8972.n49 209.834
R6810 a_n735_8972.n52 a_n735_8972.n51 209.097
R6811 a_n735_8972.n47 a_n735_8972.n0 207.859
R6812 a_n735_8972.n50 a_n735_8972.n48 207.857
R6813 a_n735_8972.n36 a_n735_8972.t50 116.401
R6814 a_n735_8972.n33 a_n735_8972.t40 116.401
R6815 a_n735_8972.n30 a_n735_8972.t44 116.401
R6816 a_n735_8972.n27 a_n735_8972.t53 116.401
R6817 a_n735_8972.n24 a_n735_8972.t41 116.401
R6818 a_n735_8972.n21 a_n735_8972.t51 116.401
R6819 a_n735_8972.n18 a_n735_8972.t45 116.401
R6820 a_n735_8972.n36 a_n735_8972.t28 115.784
R6821 a_n735_8972.n37 a_n735_8972.t47 115.784
R6822 a_n735_8972.n38 a_n735_8972.t35 115.784
R6823 a_n735_8972.n33 a_n735_8972.t46 115.784
R6824 a_n735_8972.n34 a_n735_8972.t38 115.784
R6825 a_n735_8972.n35 a_n735_8972.t27 115.784
R6826 a_n735_8972.n30 a_n735_8972.t54 115.784
R6827 a_n735_8972.n31 a_n735_8972.t42 115.784
R6828 a_n735_8972.n32 a_n735_8972.t33 115.784
R6829 a_n735_8972.n27 a_n735_8972.t31 115.784
R6830 a_n735_8972.n28 a_n735_8972.t52 115.784
R6831 a_n735_8972.n29 a_n735_8972.t37 115.784
R6832 a_n735_8972.n24 a_n735_8972.t48 115.784
R6833 a_n735_8972.n25 a_n735_8972.t39 115.784
R6834 a_n735_8972.n26 a_n735_8972.t30 115.784
R6835 a_n735_8972.n21 a_n735_8972.t49 115.784
R6836 a_n735_8972.n22 a_n735_8972.t36 115.784
R6837 a_n735_8972.n23 a_n735_8972.t32 115.784
R6838 a_n735_8972.n18 a_n735_8972.t43 115.784
R6839 a_n735_8972.n19 a_n735_8972.t34 115.784
R6840 a_n735_8972.n20 a_n735_8972.t29 115.784
R6841 a_n735_8972.n5 a_n735_8972.n4 76.6246
R6842 a_n735_8972.n11 a_n735_8972.n10 76.6229
R6843 a_n735_8972.n17 a_n735_8972.n16 76.6195
R6844 a_n735_8972.n3 a_n735_8972.n1 76.1555
R6845 a_n735_8972.n8 a_n735_8972.n6 76.1555
R6846 a_n735_8972.n14 a_n735_8972.n12 76.1555
R6847 a_n735_8972.n14 a_n735_8972.n13 75.4835
R6848 a_n735_8972.n3 a_n735_8972.n2 75.4818
R6849 a_n735_8972.n8 a_n735_8972.n7 75.4818
R6850 a_n735_8972.n49 a_n735_8972.t2 28.5655
R6851 a_n735_8972.n49 a_n735_8972.t1 28.5655
R6852 a_n735_8972.n48 a_n735_8972.t26 28.5655
R6853 a_n735_8972.n48 a_n735_8972.t24 28.5655
R6854 a_n735_8972.n0 a_n735_8972.t25 28.5655
R6855 a_n735_8972.n0 a_n735_8972.t6 28.5655
R6856 a_n735_8972.t0 a_n735_8972.n52 28.5655
R6857 a_n735_8972.n52 a_n735_8972.t5 28.5655
R6858 a_n735_8972.n45 a_n735_8972.t7 19.5762
R6859 a_n735_8972.n1 a_n735_8972.t9 17.4005
R6860 a_n735_8972.n1 a_n735_8972.t3 17.4005
R6861 a_n735_8972.n2 a_n735_8972.t4 17.4005
R6862 a_n735_8972.n2 a_n735_8972.t21 17.4005
R6863 a_n735_8972.n4 a_n735_8972.t19 17.4005
R6864 a_n735_8972.n4 a_n735_8972.t11 17.4005
R6865 a_n735_8972.n6 a_n735_8972.t15 17.4005
R6866 a_n735_8972.n6 a_n735_8972.t12 17.4005
R6867 a_n735_8972.n7 a_n735_8972.t22 17.4005
R6868 a_n735_8972.n7 a_n735_8972.t10 17.4005
R6869 a_n735_8972.n10 a_n735_8972.t13 17.4005
R6870 a_n735_8972.n10 a_n735_8972.t23 17.4005
R6871 a_n735_8972.n12 a_n735_8972.t8 17.4005
R6872 a_n735_8972.n12 a_n735_8972.t14 17.4005
R6873 a_n735_8972.n13 a_n735_8972.t17 17.4005
R6874 a_n735_8972.n13 a_n735_8972.t16 17.4005
R6875 a_n735_8972.n16 a_n735_8972.t20 17.4005
R6876 a_n735_8972.n16 a_n735_8972.t18 17.4005
R6877 a_n735_8972.n47 a_n735_8972.n46 8.00704
R6878 a_n735_8972.n45 a_n735_8972.n44 4.38516
R6879 a_n735_8972.n39 a_n735_8972.n38 3.01233
R6880 a_n735_8972.n39 a_n735_8972.n35 2.27584
R6881 a_n735_8972.n40 a_n735_8972.n32 2.27584
R6882 a_n735_8972.n41 a_n735_8972.n29 2.27584
R6883 a_n735_8972.n42 a_n735_8972.n26 2.27584
R6884 a_n735_8972.n43 a_n735_8972.n23 2.27584
R6885 a_n735_8972.n44 a_n735_8972.n20 2.27584
R6886 a_n735_8972.n46 a_n735_8972.n45 2.09073
R6887 a_n735_8972.n43 a_n735_8972.n42 1.29104
R6888 a_n735_8972.n41 a_n735_8972.n40 1.29104
R6889 a_n735_8972.n5 a_n735_8972.n3 1.07811
R6890 a_n735_8972.n9 a_n735_8972.n8 0.804722
R6891 a_n735_8972.n15 a_n735_8972.n14 0.804722
R6892 a_n735_8972.n51 a_n735_8972.n47 0.738676
R6893 a_n735_8972.n51 a_n735_8972.n50 0.736986
R6894 a_n735_8972.n38 a_n735_8972.n37 0.618487
R6895 a_n735_8972.n37 a_n735_8972.n36 0.618487
R6896 a_n735_8972.n35 a_n735_8972.n34 0.618487
R6897 a_n735_8972.n34 a_n735_8972.n33 0.618487
R6898 a_n735_8972.n32 a_n735_8972.n31 0.618487
R6899 a_n735_8972.n31 a_n735_8972.n30 0.618487
R6900 a_n735_8972.n29 a_n735_8972.n28 0.618487
R6901 a_n735_8972.n28 a_n735_8972.n27 0.618487
R6902 a_n735_8972.n26 a_n735_8972.n25 0.618487
R6903 a_n735_8972.n25 a_n735_8972.n24 0.618487
R6904 a_n735_8972.n23 a_n735_8972.n22 0.618487
R6905 a_n735_8972.n22 a_n735_8972.n21 0.618487
R6906 a_n735_8972.n20 a_n735_8972.n19 0.618487
R6907 a_n735_8972.n19 a_n735_8972.n18 0.618487
R6908 a_n735_8972.n46 a_n735_8972.n17 0.39765
R6909 a_n735_8972.n9 a_n735_8972.n5 0.27545
R6910 a_n735_8972.n17 a_n735_8972.n15 0.272317
R6911 a_n735_8972.n11 a_n735_8972.n9 0.271533
R6912 a_n735_8972.n15 a_n735_8972.n11 0.271533
R6913 a_n735_8972.n44 a_n735_8972.n43 0.182932
R6914 a_n735_8972.n42 a_n735_8972.n41 0.182932
R6915 a_n735_8972.n40 a_n735_8972.n39 0.182932
R6916 VN.n0 VN.t13 118.507
R6917 VN.n1 VN.t0 117.266
R6918 VN.n3 VN.t9 117.266
R6919 VN.n7 VN.t4 117.266
R6920 VN.n9 VN.t6 117.266
R6921 VN.n13 VN.t8 117.266
R6922 VN.n13 VN.t14 116.647
R6923 VN.n0 VN.t2 116.647
R6924 VN.n1 VN.t5 116.647
R6925 VN.n5 VN.t3 116.647
R6926 VN.n4 VN.t1 116.647
R6927 VN.n3 VN.t7 116.647
R6928 VN.n7 VN.t10 116.647
R6929 VN.n11 VN.t12 116.647
R6930 VN.n10 VN.t11 116.647
R6931 VN.n9 VN.t15 116.647
R6932 VN VN.n14 19.5341
R6933 VN.n2 VN.n0 3.8281
R6934 VN.n2 VN.n1 3.45372
R6935 VN.n8 VN.n7 3.45372
R6936 VN.n14 VN.n13 3.45372
R6937 VN.n6 VN.n5 2.21334
R6938 VN.n12 VN.n11 2.21334
R6939 VN.n4 VN.n3 1.85887
R6940 VN.n10 VN.n9 1.85887
R6941 VN.n12 VN.n8 1.00593
R6942 VN.n14 VN.n12 1.00593
R6943 VN.n6 VN.n2 0.995065
R6944 VN.n8 VN.n6 0.995065
R6945 VN.n5 VN.n4 0.618487
R6946 VN.n11 VN.n10 0.618487
R6947 a_n935_8875.n41 a_n935_8875.n35 203.368
R6948 a_n935_8875.n6 a_n935_8875.n4 203.368
R6949 a_n935_8875.n19 a_n935_8875.n13 203.368
R6950 a_n935_8875.n27 a_n935_8875.n25 203.368
R6951 a_n935_8875.n15 a_n935_8875.t36 116.401
R6952 a_n935_8875.n37 a_n935_8875.t35 116.401
R6953 a_n935_8875.n11 a_n935_8875.t39 115.784
R6954 a_n935_8875.n10 a_n935_8875.t40 115.784
R6955 a_n935_8875.n15 a_n935_8875.t34 115.784
R6956 a_n935_8875.n32 a_n935_8875.t37 115.784
R6957 a_n935_8875.n31 a_n935_8875.t38 115.784
R6958 a_n935_8875.n37 a_n935_8875.t41 115.784
R6959 a_n935_8875.n5 a_n935_8875.t20 113.578
R6960 a_n935_8875.n26 a_n935_8875.t22 113.578
R6961 a_n935_8875.n8 a_n935_8875.t24 113.532
R6962 a_n935_8875.n21 a_n935_8875.t28 113.532
R6963 a_n935_8875.n14 a_n935_8875.t26 113.532
R6964 a_n935_8875.n29 a_n935_8875.t30 113.532
R6965 a_n935_8875.n43 a_n935_8875.t32 113.532
R6966 a_n935_8875.n36 a_n935_8875.t18 113.532
R6967 a_n935_8875.n55 a_n935_8875.n54 76.6009
R6968 a_n935_8875.n59 a_n935_8875.n58 76.3312
R6969 a_n935_8875.n56 a_n935_8875.n50 76.3312
R6970 a_n935_8875.n53 a_n935_8875.n51 76.1487
R6971 a_n935_8875.n49 a_n935_8875.n47 76.1487
R6972 a_n935_8875.n2 a_n935_8875.n0 76.1487
R6973 a_n935_8875.n53 a_n935_8875.n52 75.4751
R6974 a_n935_8875.n49 a_n935_8875.n48 75.4751
R6975 a_n935_8875.n2 a_n935_8875.n1 75.4751
R6976 a_n935_8875.n4 a_n935_8875.t21 28.5655
R6977 a_n935_8875.n4 a_n935_8875.t25 28.5655
R6978 a_n935_8875.n13 a_n935_8875.t27 28.5655
R6979 a_n935_8875.n13 a_n935_8875.t29 28.5655
R6980 a_n935_8875.n25 a_n935_8875.t23 28.5655
R6981 a_n935_8875.n25 a_n935_8875.t31 28.5655
R6982 a_n935_8875.n35 a_n935_8875.t19 28.5655
R6983 a_n935_8875.n35 a_n935_8875.t33 28.5655
R6984 a_n935_8875.n54 a_n935_8875.t7 17.4005
R6985 a_n935_8875.n54 a_n935_8875.t1 17.4005
R6986 a_n935_8875.n52 a_n935_8875.t4 17.4005
R6987 a_n935_8875.n52 a_n935_8875.t3 17.4005
R6988 a_n935_8875.n51 a_n935_8875.t9 17.4005
R6989 a_n935_8875.n51 a_n935_8875.t0 17.4005
R6990 a_n935_8875.n50 a_n935_8875.t11 17.4005
R6991 a_n935_8875.n50 a_n935_8875.t5 17.4005
R6992 a_n935_8875.n48 a_n935_8875.t14 17.4005
R6993 a_n935_8875.n48 a_n935_8875.t12 17.4005
R6994 a_n935_8875.n47 a_n935_8875.t6 17.4005
R6995 a_n935_8875.n47 a_n935_8875.t8 17.4005
R6996 a_n935_8875.n1 a_n935_8875.t13 17.4005
R6997 a_n935_8875.n1 a_n935_8875.t16 17.4005
R6998 a_n935_8875.n0 a_n935_8875.t17 17.4005
R6999 a_n935_8875.n0 a_n935_8875.t2 17.4005
R7000 a_n935_8875.t15 a_n935_8875.n59 17.4005
R7001 a_n935_8875.n59 a_n935_8875.t10 17.4005
R7002 a_n935_8875.n46 a_n935_8875.n45 12.8828
R7003 a_n935_8875.n9 a_n935_8875.n8 4.5872
R7004 a_n935_8875.n22 a_n935_8875.n21 4.5872
R7005 a_n935_8875.n16 a_n935_8875.n14 4.5872
R7006 a_n935_8875.n30 a_n935_8875.n29 4.5872
R7007 a_n935_8875.n44 a_n935_8875.n43 4.5872
R7008 a_n935_8875.n38 a_n935_8875.n36 4.5872
R7009 a_n935_8875.n7 a_n935_8875.n3 4.5005
R7010 a_n935_8875.n18 a_n935_8875.n17 4.5005
R7011 a_n935_8875.n20 a_n935_8875.n12 4.5005
R7012 a_n935_8875.n28 a_n935_8875.n24 4.5005
R7013 a_n935_8875.n42 a_n935_8875.n34 4.5005
R7014 a_n935_8875.n40 a_n935_8875.n39 4.5005
R7015 a_n935_8875.n5 a_n935_8875.n3 2.73978
R7016 a_n935_8875.n26 a_n935_8875.n24 2.73978
R7017 a_n935_8875.n23 a_n935_8875.n11 2.44892
R7018 a_n935_8875.n33 a_n935_8875.n32 2.3143
R7019 a_n935_8875.n23 a_n935_8875.n22 2.22887
R7020 a_n935_8875.n45 a_n935_8875.n44 2.22887
R7021 a_n935_8875.n33 a_n935_8875.n23 1.71204
R7022 a_n935_8875.n11 a_n935_8875.n10 0.618487
R7023 a_n935_8875.n32 a_n935_8875.n31 0.618487
R7024 a_n935_8875.n10 a_n935_8875.n9 0.533051
R7025 a_n935_8875.n16 a_n935_8875.n15 0.533051
R7026 a_n935_8875.n31 a_n935_8875.n30 0.533051
R7027 a_n935_8875.n38 a_n935_8875.n37 0.533051
R7028 a_n935_8875.n55 a_n935_8875.n53 0.521417
R7029 a_n935_8875.n57 a_n935_8875.n49 0.521417
R7030 a_n935_8875.n46 a_n935_8875.n2 0.521417
R7031 a_n935_8875.n17 a_n935_8875.n12 0.447615
R7032 a_n935_8875.n39 a_n935_8875.n34 0.447615
R7033 a_n935_8875.n56 a_n935_8875.n55 0.269162
R7034 a_n935_8875.n6 a_n935_8875.n5 0.2663
R7035 a_n935_8875.n27 a_n935_8875.n26 0.2663
R7036 a_n935_8875.n58 a_n935_8875.n46 0.265986
R7037 a_n935_8875.n58 a_n935_8875.n57 0.265986
R7038 a_n935_8875.n57 a_n935_8875.n56 0.265986
R7039 a_n935_8875.n7 a_n935_8875.n6 0.224058
R7040 a_n935_8875.n19 a_n935_8875.n18 0.224058
R7041 a_n935_8875.n20 a_n935_8875.n19 0.224058
R7042 a_n935_8875.n28 a_n935_8875.n27 0.224058
R7043 a_n935_8875.n41 a_n935_8875.n40 0.224058
R7044 a_n935_8875.n42 a_n935_8875.n41 0.224058
R7045 a_n935_8875.n9 a_n935_8875.n3 0.173577
R7046 a_n935_8875.n17 a_n935_8875.n16 0.173577
R7047 a_n935_8875.n22 a_n935_8875.n12 0.173577
R7048 a_n935_8875.n30 a_n935_8875.n24 0.173577
R7049 a_n935_8875.n39 a_n935_8875.n38 0.173577
R7050 a_n935_8875.n44 a_n935_8875.n34 0.173577
R7051 a_n935_8875.n45 a_n935_8875.n33 0.135115
R7052 a_n935_8875.n8 a_n935_8875.n7 0.0871986
R7053 a_n935_8875.n18 a_n935_8875.n14 0.0871986
R7054 a_n935_8875.n21 a_n935_8875.n20 0.0871986
R7055 a_n935_8875.n29 a_n935_8875.n28 0.0871986
R7056 a_n935_8875.n40 a_n935_8875.n36 0.0871986
R7057 a_n935_8875.n43 a_n935_8875.n42 0.0871986
R7058 a_9909_7861.t0 a_9909_7861.t1 21.0809
C0 IBIAS VDD 0.01133f
C1 IBIAS VN 0.30289f
C2 EN VDD 0.03838f
C3 EN VN 0.10946f
C4 EN VP 0.15973f
C5 IBIAS VOUT 10.8674f
C6 EN VOUT 3.59173f
C7 IBIAS EN 49.9753f
C8 VDD VN 0.12959f
C9 VDD VP 0.88136f
C10 VN VP 8.1017f
C11 VDD VOUT 3.03127f
C12 EN VSS 58.70063f
C13 IBIAS VSS 63.26237f
C14 VOUT VSS 74.14656f
C15 VP VSS 13.6618f
C16 VN VSS 11.84216f
C17 VDD VSS 41.71331f
C18 a_9909_7861.t1 VSS 0.22264p
C19 a_9909_7861.t0 VSS 0.75527f
C20 a_n935_8875.t17 VSS 0.0162f
C21 a_n935_8875.t2 VSS 0.0162f
C22 a_n935_8875.n0 VSS 0.05074f
C23 a_n935_8875.t13 VSS 0.0162f
C24 a_n935_8875.t16 VSS 0.0162f
C25 a_n935_8875.n1 VSS 0.04731f
C26 a_n935_8875.n2 VSS 0.91776f
C27 a_n935_8875.n3 VSS 0.0928f
C28 a_n935_8875.t21 VSS 0.0162f
C29 a_n935_8875.t25 VSS 0.0162f
C30 a_n935_8875.n4 VSS 0.0339f
C31 a_n935_8875.t20 VSS 0.18352f
C32 a_n935_8875.n5 VSS 0.12983f
C33 a_n935_8875.n6 VSS 0.14005f
C34 a_n935_8875.n7 VSS 0.03712f
C35 a_n935_8875.t24 VSS 0.18349f
C36 a_n935_8875.n8 VSS 0.08677f
C37 a_n935_8875.n9 VSS 0.04427f
C38 a_n935_8875.t40 VSS 0.18586f
C39 a_n935_8875.n10 VSS 0.18972f
C40 a_n935_8875.t39 VSS 0.18586f
C41 a_n935_8875.n11 VSS 0.30068f
C42 a_n935_8875.n12 VSS 0.03747f
C43 a_n935_8875.t27 VSS 0.0162f
C44 a_n935_8875.t29 VSS 0.0162f
C45 a_n935_8875.n13 VSS 0.0339f
C46 a_n935_8875.t26 VSS 0.18349f
C47 a_n935_8875.n14 VSS 0.08677f
C48 a_n935_8875.t36 VSS 0.18686f
C49 a_n935_8875.t34 VSS 0.18586f
C50 a_n935_8875.n15 VSS 0.37614f
C51 a_n935_8875.n16 VSS 0.04427f
C52 a_n935_8875.n17 VSS 0.03747f
C53 a_n935_8875.n18 VSS 0.03712f
C54 a_n935_8875.n19 VSS 0.13415f
C55 a_n935_8875.n20 VSS 0.03712f
C56 a_n935_8875.t28 VSS 0.18349f
C57 a_n935_8875.n21 VSS 0.08677f
C58 a_n935_8875.n22 VSS 0.14577f
C59 a_n935_8875.n23 VSS 0.29849f
C60 a_n935_8875.n24 VSS 0.0928f
C61 a_n935_8875.t23 VSS 0.0162f
C62 a_n935_8875.t31 VSS 0.0162f
C63 a_n935_8875.n25 VSS 0.0339f
C64 a_n935_8875.t22 VSS 0.18352f
C65 a_n935_8875.n26 VSS 0.12983f
C66 a_n935_8875.n27 VSS 0.14005f
C67 a_n935_8875.n28 VSS 0.03712f
C68 a_n935_8875.t30 VSS 0.18349f
C69 a_n935_8875.n29 VSS 0.08677f
C70 a_n935_8875.n30 VSS 0.04427f
C71 a_n935_8875.t38 VSS 0.18586f
C72 a_n935_8875.n31 VSS 0.18972f
C73 a_n935_8875.t37 VSS 0.18586f
C74 a_n935_8875.n32 VSS 0.29808f
C75 a_n935_8875.n33 VSS 0.25912f
C76 a_n935_8875.n34 VSS 0.03747f
C77 a_n935_8875.t19 VSS 0.0162f
C78 a_n935_8875.t33 VSS 0.0162f
C79 a_n935_8875.n35 VSS 0.0339f
C80 a_n935_8875.t18 VSS 0.18349f
C81 a_n935_8875.n36 VSS 0.08677f
C82 a_n935_8875.t35 VSS 0.18686f
C83 a_n935_8875.t41 VSS 0.18586f
C84 a_n935_8875.n37 VSS 0.37614f
C85 a_n935_8875.n38 VSS 0.04427f
C86 a_n935_8875.n39 VSS 0.03747f
C87 a_n935_8875.n40 VSS 0.03712f
C88 a_n935_8875.n41 VSS 0.13415f
C89 a_n935_8875.n42 VSS 0.03712f
C90 a_n935_8875.t32 VSS 0.18349f
C91 a_n935_8875.n43 VSS 0.08677f
C92 a_n935_8875.n44 VSS 0.14577f
C93 a_n935_8875.n45 VSS 1.43716f
C94 a_n935_8875.n46 VSS 1.14056f
C95 a_n935_8875.t6 VSS 0.0162f
C96 a_n935_8875.t8 VSS 0.0162f
C97 a_n935_8875.n47 VSS 0.05083f
C98 a_n935_8875.t14 VSS 0.0162f
C99 a_n935_8875.t12 VSS 0.0162f
C100 a_n935_8875.n48 VSS 0.04731f
C101 a_n935_8875.n49 VSS 0.91932f
C102 a_n935_8875.t11 VSS 0.0162f
C103 a_n935_8875.t5 VSS 0.0162f
C104 a_n935_8875.n50 VSS 0.0523f
C105 a_n935_8875.t9 VSS 0.0162f
C106 a_n935_8875.t0 VSS 0.0162f
C107 a_n935_8875.n51 VSS 0.05074f
C108 a_n935_8875.t4 VSS 0.0162f
C109 a_n935_8875.t3 VSS 0.0162f
C110 a_n935_8875.n52 VSS 0.04731f
C111 a_n935_8875.n53 VSS 0.91776f
C112 a_n935_8875.t7 VSS 0.0162f
C113 a_n935_8875.t1 VSS 0.0162f
C114 a_n935_8875.n54 VSS 0.05493f
C115 a_n935_8875.n55 VSS 1.03058f
C116 a_n935_8875.n56 VSS 0.8237f
C117 a_n935_8875.n57 VSS 0.27938f
C118 a_n935_8875.n58 VSS 0.82267f
C119 a_n935_8875.t10 VSS 0.0162f
C120 a_n935_8875.n59 VSS 0.0523f
C121 a_n935_8875.t15 VSS 0.0162f
C122 VN.t13 VSS 0.24256f
C123 VN.t2 VSS 0.23725f
C124 VN.n0 VSS 0.92639f
C125 VN.t0 VSS 0.23838f
C126 VN.t5 VSS 0.23712f
C127 VN.n1 VSS 0.70238f
C128 VN.n2 VSS 0.59951f
C129 VN.t9 VSS 0.23838f
C130 VN.t7 VSS 0.23712f
C131 VN.n3 VSS 0.58122f
C132 VN.t1 VSS 0.23712f
C133 VN.n4 VSS 0.34446f
C134 VN.t3 VSS 0.23712f
C135 VN.n5 VSS 0.37114f
C136 VN.n6 VSS 0.29549f
C137 VN.t4 VSS 0.23838f
C138 VN.t10 VSS 0.23712f
C139 VN.n7 VSS 0.70238f
C140 VN.n8 VSS 0.3904f
C141 VN.t6 VSS 0.23838f
C142 VN.t15 VSS 0.23712f
C143 VN.n9 VSS 0.58122f
C144 VN.t11 VSS 0.23712f
C145 VN.n10 VSS 0.34446f
C146 VN.t12 VSS 0.23712f
C147 VN.n11 VSS 0.37114f
C148 VN.n12 VSS 0.29678f
C149 VN.t8 VSS 0.23838f
C150 VN.t14 VSS 0.23712f
C151 VN.n13 VSS 0.70238f
C152 VN.n14 VSS 1.48757f
C153 a_n735_8972.t25 VSS 0.01366f
C154 a_n735_8972.t6 VSS 0.01366f
C155 a_n735_8972.n0 VSS 0.03271f
C156 a_n735_8972.t9 VSS 0.01366f
C157 a_n735_8972.t3 VSS 0.01366f
C158 a_n735_8972.n1 VSS 0.04286f
C159 a_n735_8972.t4 VSS 0.01366f
C160 a_n735_8972.t21 VSS 0.01366f
C161 a_n735_8972.n2 VSS 0.03996f
C162 a_n735_8972.n3 VSS 0.91801f
C163 a_n735_8972.t19 VSS 0.01366f
C164 a_n735_8972.t11 VSS 0.01366f
C165 a_n735_8972.n4 VSS 0.04666f
C166 a_n735_8972.n5 VSS 1.04866f
C167 a_n735_8972.t15 VSS 0.01366f
C168 a_n735_8972.t12 VSS 0.01366f
C169 a_n735_8972.n6 VSS 0.04286f
C170 a_n735_8972.t22 VSS 0.01366f
C171 a_n735_8972.t10 VSS 0.01366f
C172 a_n735_8972.n7 VSS 0.03996f
C173 a_n735_8972.n8 VSS 0.84993f
C174 a_n735_8972.n9 VSS 0.31753f
C175 a_n735_8972.t13 VSS 0.01366f
C176 a_n735_8972.t23 VSS 0.01366f
C177 a_n735_8972.n10 VSS 0.04665f
C178 a_n735_8972.n11 VSS 0.84725f
C179 a_n735_8972.t8 VSS 0.01366f
C180 a_n735_8972.t14 VSS 0.01366f
C181 a_n735_8972.n12 VSS 0.04286f
C182 a_n735_8972.t17 VSS 0.01366f
C183 a_n735_8972.t16 VSS 0.01366f
C184 a_n735_8972.n13 VSS 0.03996f
C185 a_n735_8972.n14 VSS 0.84993f
C186 a_n735_8972.n15 VSS 0.31696f
C187 a_n735_8972.t20 VSS 0.01366f
C188 a_n735_8972.t18 VSS 0.01366f
C189 a_n735_8972.n16 VSS 0.04665f
C190 a_n735_8972.n17 VSS 0.87015f
C191 a_n735_8972.t7 VSS 0.89417f
C192 a_n735_8972.t45 VSS 0.1575f
C193 a_n735_8972.t43 VSS 0.15669f
C194 a_n735_8972.n18 VSS 0.3169f
C195 a_n735_8972.t34 VSS 0.15669f
C196 a_n735_8972.n19 VSS 0.1651f
C197 a_n735_8972.t29 VSS 0.15669f
C198 a_n735_8972.n20 VSS 0.24934f
C199 a_n735_8972.t51 VSS 0.1575f
C200 a_n735_8972.t49 VSS 0.15669f
C201 a_n735_8972.n21 VSS 0.3169f
C202 a_n735_8972.t36 VSS 0.15669f
C203 a_n735_8972.n22 VSS 0.1651f
C204 a_n735_8972.t32 VSS 0.15669f
C205 a_n735_8972.n23 VSS 0.24934f
C206 a_n735_8972.t41 VSS 0.1575f
C207 a_n735_8972.t48 VSS 0.15669f
C208 a_n735_8972.n24 VSS 0.3169f
C209 a_n735_8972.t39 VSS 0.15669f
C210 a_n735_8972.n25 VSS 0.1651f
C211 a_n735_8972.t30 VSS 0.15669f
C212 a_n735_8972.n26 VSS 0.24934f
C213 a_n735_8972.t53 VSS 0.1575f
C214 a_n735_8972.t31 VSS 0.15669f
C215 a_n735_8972.n27 VSS 0.3169f
C216 a_n735_8972.t52 VSS 0.15669f
C217 a_n735_8972.n28 VSS 0.1651f
C218 a_n735_8972.t37 VSS 0.15669f
C219 a_n735_8972.n29 VSS 0.24934f
C220 a_n735_8972.t44 VSS 0.1575f
C221 a_n735_8972.t54 VSS 0.15669f
C222 a_n735_8972.n30 VSS 0.3169f
C223 a_n735_8972.t42 VSS 0.15669f
C224 a_n735_8972.n31 VSS 0.1651f
C225 a_n735_8972.t33 VSS 0.15669f
C226 a_n735_8972.n32 VSS 0.24934f
C227 a_n735_8972.t40 VSS 0.1575f
C228 a_n735_8972.t46 VSS 0.15669f
C229 a_n735_8972.n33 VSS 0.3169f
C230 a_n735_8972.t38 VSS 0.15669f
C231 a_n735_8972.n34 VSS 0.1651f
C232 a_n735_8972.t27 VSS 0.15669f
C233 a_n735_8972.n35 VSS 0.24934f
C234 a_n735_8972.t50 VSS 0.1575f
C235 a_n735_8972.t28 VSS 0.15669f
C236 a_n735_8972.n36 VSS 0.3169f
C237 a_n735_8972.t47 VSS 0.15669f
C238 a_n735_8972.n37 VSS 0.1651f
C239 a_n735_8972.t35 VSS 0.15669f
C240 a_n735_8972.n38 VSS 0.32068f
C241 a_n735_8972.n39 VSS 0.43128f
C242 a_n735_8972.n40 VSS 0.26804f
C243 a_n735_8972.n41 VSS 0.26804f
C244 a_n735_8972.n42 VSS 0.26804f
C245 a_n735_8972.n43 VSS 0.26804f
C246 a_n735_8972.n44 VSS 0.32368f
C247 a_n735_8972.n45 VSS 1.79294f
C248 a_n735_8972.n46 VSS 1.73175f
C249 a_n735_8972.n47 VSS 0.86736f
C250 a_n735_8972.t26 VSS 0.01366f
C251 a_n735_8972.t24 VSS 0.01366f
C252 a_n735_8972.n48 VSS 0.03271f
C253 a_n735_8972.t2 VSS 0.01366f
C254 a_n735_8972.t1 VSS 0.01366f
C255 a_n735_8972.n49 VSS 0.03783f
C256 a_n735_8972.n50 VSS 1.22547f
C257 a_n735_8972.n51 VSS 0.67677f
C258 a_n735_8972.t5 VSS 0.01366f
C259 a_n735_8972.n52 VSS 0.03547f
C260 a_n735_8972.t0 VSS 0.01366f
C261 VP.t14 VSS 0.23122f
C262 VP.t2 VSS 0.22624f
C263 VP.n0 VSS 0.86272f
C264 VP.t12 VSS 0.22744f
C265 VP.t4 VSS 0.22624f
C266 VP.n1 VSS 0.66072f
C267 VP.n2 VSS 0.55267f
C268 VP.t11 VSS 0.22744f
C269 VP.t8 VSS 0.22624f
C270 VP.n3 VSS 0.55455f
C271 VP.t13 VSS 0.22624f
C272 VP.n4 VSS 0.32865f
C273 VP.t1 VSS 0.22624f
C274 VP.n5 VSS 0.34467f
C275 VP.n6 VSS 0.27314f
C276 VP.t0 VSS 0.22743f
C277 VP.t10 VSS 0.22624f
C278 VP.n7 VSS 0.65941f
C279 VP.n8 VSS 0.36245f
C280 VP.t9 VSS 0.22744f
C281 VP.t15 VSS 0.22624f
C282 VP.n9 VSS 0.55455f
C283 VP.t7 VSS 0.22624f
C284 VP.n10 VSS 0.32865f
C285 VP.t6 VSS 0.22624f
C286 VP.n11 VSS 0.34467f
C287 VP.n12 VSS 0.27252f
C288 VP.t5 VSS 0.22744f
C289 VP.t3 VSS 0.22624f
C290 VP.n13 VSS 0.66072f
C291 VP.n14 VSS 1.99935f
C292 a_n1962_4406.t89 VSS 0.02309f
C293 a_n1962_4406.t22 VSS 0.02309f
C294 a_n1962_4406.t3 VSS 0.02309f
C295 a_n1962_4406.n0 VSS 0.05448f
C296 a_n1962_4406.t115 VSS 0.02309f
C297 a_n1962_4406.t30 VSS 0.02309f
C298 a_n1962_4406.n1 VSS 0.05185f
C299 a_n1962_4406.n2 VSS 0.31248f
C300 a_n1962_4406.t54 VSS 0.02309f
C301 a_n1962_4406.t57 VSS 0.02309f
C302 a_n1962_4406.n3 VSS 0.05448f
C303 a_n1962_4406.t25 VSS 0.02309f
C304 a_n1962_4406.t96 VSS 0.02309f
C305 a_n1962_4406.n4 VSS 0.05185f
C306 a_n1962_4406.n5 VSS 0.31248f
C307 a_n1962_4406.t31 VSS 0.02309f
C308 a_n1962_4406.t33 VSS 0.02309f
C309 a_n1962_4406.n6 VSS 0.05448f
C310 a_n1962_4406.t90 VSS 0.02309f
C311 a_n1962_4406.t15 VSS 0.02309f
C312 a_n1962_4406.n7 VSS 0.05185f
C313 a_n1962_4406.n8 VSS 0.36496f
C314 a_n1962_4406.t48 VSS 0.02309f
C315 a_n1962_4406.t116 VSS 0.02309f
C316 a_n1962_4406.n9 VSS 0.05185f
C317 a_n1962_4406.n10 VSS 0.20376f
C318 a_n1962_4406.t91 VSS 0.02309f
C319 a_n1962_4406.t16 VSS 0.02309f
C320 a_n1962_4406.n11 VSS 0.05185f
C321 a_n1962_4406.n12 VSS 0.20376f
C322 a_n1962_4406.t49 VSS 0.02309f
C323 a_n1962_4406.t117 VSS 0.02309f
C324 a_n1962_4406.n13 VSS 0.05185f
C325 a_n1962_4406.n14 VSS 0.20376f
C326 a_n1962_4406.t103 VSS 0.02309f
C327 a_n1962_4406.t37 VSS 0.02309f
C328 a_n1962_4406.n15 VSS 0.05185f
C329 a_n1962_4406.n16 VSS 0.20376f
C330 a_n1962_4406.t10 VSS 0.02309f
C331 a_n1962_4406.t86 VSS 0.02309f
C332 a_n1962_4406.n17 VSS 0.05185f
C333 a_n1962_4406.n18 VSS 0.15234f
C334 a_n1962_4406.t42 VSS 0.02309f
C335 a_n1962_4406.t79 VSS 0.02309f
C336 a_n1962_4406.n19 VSS 0.05448f
C337 a_n1962_4406.t87 VSS 0.02309f
C338 a_n1962_4406.t27 VSS 0.02309f
C339 a_n1962_4406.n20 VSS 0.05185f
C340 a_n1962_4406.n21 VSS 0.31291f
C341 a_n1962_4406.t12 VSS 0.02309f
C342 a_n1962_4406.t66 VSS 0.02309f
C343 a_n1962_4406.n22 VSS 0.05255f
C344 a_n1962_4406.t23 VSS 0.02309f
C345 a_n1962_4406.t68 VSS 0.02309f
C346 a_n1962_4406.n23 VSS 0.05448f
C347 a_n1962_4406.t81 VSS 0.02309f
C348 a_n1962_4406.t6 VSS 0.02309f
C349 a_n1962_4406.n24 VSS 0.05185f
C350 a_n1962_4406.n25 VSS 0.36496f
C351 a_n1962_4406.t34 VSS 0.02309f
C352 a_n1962_4406.t107 VSS 0.02309f
C353 a_n1962_4406.n26 VSS 0.05185f
C354 a_n1962_4406.n27 VSS 0.20376f
C355 a_n1962_4406.t82 VSS 0.02309f
C356 a_n1962_4406.t7 VSS 0.02309f
C357 a_n1962_4406.n28 VSS 0.05185f
C358 a_n1962_4406.n29 VSS 0.20376f
C359 a_n1962_4406.t35 VSS 0.02309f
C360 a_n1962_4406.t108 VSS 0.02309f
C361 a_n1962_4406.n30 VSS 0.05185f
C362 a_n1962_4406.n31 VSS 0.20376f
C363 a_n1962_4406.t94 VSS 0.02309f
C364 a_n1962_4406.t28 VSS 0.02309f
C365 a_n1962_4406.n32 VSS 0.05185f
C366 a_n1962_4406.n33 VSS 0.20376f
C367 a_n1962_4406.t55 VSS 0.02309f
C368 a_n1962_4406.t122 VSS 0.02309f
C369 a_n1962_4406.n34 VSS 0.05185f
C370 a_n1962_4406.n35 VSS 0.15465f
C371 a_n1962_4406.t44 VSS 0.02309f
C372 a_n1962_4406.t65 VSS 0.02309f
C373 a_n1962_4406.n36 VSS 0.05299f
C374 a_n1962_4406.t8 VSS 0.02309f
C375 a_n1962_4406.t72 VSS 0.02309f
C376 a_n1962_4406.n37 VSS 0.05494f
C377 a_n1962_4406.t109 VSS 0.02309f
C378 a_n1962_4406.t61 VSS 0.02309f
C379 a_n1962_4406.n38 VSS 0.05185f
C380 a_n1962_4406.n39 VSS 0.39307f
C381 a_n1962_4406.t9 VSS 0.02309f
C382 a_n1962_4406.t73 VSS 0.02309f
C383 a_n1962_4406.n40 VSS 0.05185f
C384 a_n1962_4406.n41 VSS 0.20376f
C385 a_n1962_4406.t110 VSS 0.02309f
C386 a_n1962_4406.t62 VSS 0.02309f
C387 a_n1962_4406.n42 VSS 0.05185f
C388 a_n1962_4406.n43 VSS 0.20376f
C389 a_n1962_4406.t29 VSS 0.02309f
C390 a_n1962_4406.t77 VSS 0.02309f
C391 a_n1962_4406.n44 VSS 0.05185f
C392 a_n1962_4406.n45 VSS 0.20376f
C393 a_n1962_4406.t123 VSS 0.02309f
C394 a_n1962_4406.t69 VSS 0.02309f
C395 a_n1962_4406.n46 VSS 0.05185f
C396 a_n1962_4406.n47 VSS 0.15465f
C397 a_n1962_4406.n48 VSS 0.32645f
C398 a_n1962_4406.n49 VSS 0.17936f
C399 a_n1962_4406.t111 VSS 0.02309f
C400 a_n1962_4406.t43 VSS 0.02309f
C401 a_n1962_4406.n50 VSS 0.05185f
C402 a_n1962_4406.n51 VSS 0.11823f
C403 a_n1962_4406.n52 VSS 0.29057f
C404 a_n1962_4406.n53 VSS 0.17949f
C405 a_n1962_4406.t41 VSS 0.02309f
C406 a_n1962_4406.t120 VSS 0.02309f
C407 a_n1962_4406.n54 VSS 0.05185f
C408 a_n1962_4406.n55 VSS 0.12045f
C409 a_n1962_4406.t24 VSS 0.02309f
C410 a_n1962_4406.t32 VSS 0.02309f
C411 a_n1962_4406.n56 VSS 0.05448f
C412 a_n1962_4406.t4 VSS 0.02309f
C413 a_n1962_4406.t92 VSS 0.02309f
C414 a_n1962_4406.n57 VSS 0.05185f
C415 a_n1962_4406.n58 VSS 0.36496f
C416 a_n1962_4406.t104 VSS 0.02309f
C417 a_n1962_4406.t50 VSS 0.02309f
C418 a_n1962_4406.n59 VSS 0.05185f
C419 a_n1962_4406.n60 VSS 0.20376f
C420 a_n1962_4406.t5 VSS 0.02309f
C421 a_n1962_4406.t93 VSS 0.02309f
C422 a_n1962_4406.n61 VSS 0.05185f
C423 a_n1962_4406.n62 VSS 0.20376f
C424 a_n1962_4406.t105 VSS 0.02309f
C425 a_n1962_4406.t51 VSS 0.02309f
C426 a_n1962_4406.n63 VSS 0.05185f
C427 a_n1962_4406.n64 VSS 0.20376f
C428 a_n1962_4406.t26 VSS 0.02309f
C429 a_n1962_4406.t106 VSS 0.02309f
C430 a_n1962_4406.n65 VSS 0.05185f
C431 a_n1962_4406.n66 VSS 0.20376f
C432 a_n1962_4406.t121 VSS 0.02309f
C433 a_n1962_4406.t11 VSS 0.02309f
C434 a_n1962_4406.n67 VSS 0.05185f
C435 a_n1962_4406.n68 VSS 0.15234f
C436 a_n1962_4406.n69 VSS 0.17945f
C437 a_n1962_4406.n70 VSS 0.17945f
C438 a_n1962_4406.t119 VSS 0.02309f
C439 a_n1962_4406.t56 VSS 0.02309f
C440 a_n1962_4406.n71 VSS 0.05185f
C441 a_n1962_4406.n72 VSS 0.12085f
C442 a_n1962_4406.n73 VSS 0.17952f
C443 a_n1962_4406.n74 VSS 0.17952f
C444 a_n1962_4406.t20 VSS 0.02309f
C445 a_n1962_4406.t80 VSS 0.02309f
C446 a_n1962_4406.n75 VSS 0.05185f
C447 a_n1962_4406.n76 VSS 0.12185f
C448 a_n1962_4406.t70 VSS 0.02309f
C449 a_n1962_4406.t39 VSS 0.02309f
C450 a_n1962_4406.n77 VSS 0.05448f
C451 a_n1962_4406.t52 VSS 0.02309f
C452 a_n1962_4406.t84 VSS 0.02309f
C453 a_n1962_4406.n78 VSS 0.05185f
C454 a_n1962_4406.n79 VSS 0.3114f
C455 a_n1962_4406.t75 VSS 0.02309f
C456 a_n1962_4406.t53 VSS 0.02309f
C457 a_n1962_4406.n80 VSS 0.05268f
C458 a_n1962_4406.t63 VSS 0.02309f
C459 a_n1962_4406.t19 VSS 0.02309f
C460 a_n1962_4406.n81 VSS 0.05494f
C461 a_n1962_4406.t74 VSS 0.02309f
C462 a_n1962_4406.t114 VSS 0.02309f
C463 a_n1962_4406.n82 VSS 0.05185f
C464 a_n1962_4406.n83 VSS 0.39307f
C465 a_n1962_4406.t64 VSS 0.02309f
C466 a_n1962_4406.t21 VSS 0.02309f
C467 a_n1962_4406.n84 VSS 0.05185f
C468 a_n1962_4406.n85 VSS 0.20376f
C469 a_n1962_4406.t78 VSS 0.02309f
C470 a_n1962_4406.t85 VSS 0.02309f
C471 a_n1962_4406.n86 VSS 0.05185f
C472 a_n1962_4406.n87 VSS 0.20376f
C473 a_n1962_4406.t71 VSS 0.02309f
C474 a_n1962_4406.t40 VSS 0.02309f
C475 a_n1962_4406.n88 VSS 0.05185f
C476 a_n1962_4406.n89 VSS 0.20376f
C477 a_n1962_4406.t67 VSS 0.02309f
C478 a_n1962_4406.t97 VSS 0.02309f
C479 a_n1962_4406.n90 VSS 0.05185f
C480 a_n1962_4406.n91 VSS 0.1638f
C481 a_n1962_4406.n92 VSS 0.31762f
C482 a_n1962_4406.n93 VSS 0.17959f
C483 a_n1962_4406.t95 VSS 0.02309f
C484 a_n1962_4406.t36 VSS 0.02309f
C485 a_n1962_4406.n94 VSS 0.05185f
C486 a_n1962_4406.n95 VSS 0.12285f
C487 a_n1962_4406.t76 VSS 0.02309f
C488 a_n1962_4406.t0 VSS 0.02309f
C489 a_n1962_4406.n96 VSS 0.05449f
C490 a_n1962_4406.t14 VSS 0.02309f
C491 a_n1962_4406.t100 VSS 0.02309f
C492 a_n1962_4406.n97 VSS 0.05185f
C493 a_n1962_4406.n98 VSS 0.36532f
C494 a_n1962_4406.t113 VSS 0.02309f
C495 a_n1962_4406.t1 VSS 0.02309f
C496 a_n1962_4406.n99 VSS 0.05185f
C497 a_n1962_4406.n100 VSS 0.20376f
C498 a_n1962_4406.t17 VSS 0.02309f
C499 a_n1962_4406.t101 VSS 0.02309f
C500 a_n1962_4406.n101 VSS 0.05185f
C501 a_n1962_4406.n102 VSS 0.20376f
C502 a_n1962_4406.t83 VSS 0.02309f
C503 a_n1962_4406.t18 VSS 0.02309f
C504 a_n1962_4406.n103 VSS 0.05185f
C505 a_n1962_4406.n104 VSS 0.20376f
C506 a_n1962_4406.t38 VSS 0.02309f
C507 a_n1962_4406.t118 VSS 0.02309f
C508 a_n1962_4406.n105 VSS 0.05185f
C509 a_n1962_4406.n106 VSS 0.15127f
C510 a_n1962_4406.n107 VSS 0.17952f
C511 a_n1962_4406.n108 VSS 0.17952f
C512 a_n1962_4406.t102 VSS 0.02309f
C513 a_n1962_4406.t13 VSS 0.02309f
C514 a_n1962_4406.n109 VSS 0.05185f
C515 a_n1962_4406.n110 VSS 0.15127f
C516 a_n1962_4406.t2 VSS 0.02309f
C517 a_n1962_4406.t112 VSS 0.02309f
C518 a_n1962_4406.n111 VSS 0.05185f
C519 a_n1962_4406.n112 VSS 0.20376f
C520 a_n1962_4406.t60 VSS 0.02309f
C521 a_n1962_4406.t45 VSS 0.02309f
C522 a_n1962_4406.n113 VSS 0.05448f
C523 a_n1962_4406.t46 VSS 0.02309f
C524 a_n1962_4406.t98 VSS 0.02309f
C525 a_n1962_4406.n114 VSS 0.05185f
C526 a_n1962_4406.n115 VSS 0.36496f
C527 a_n1962_4406.t88 VSS 0.02309f
C528 a_n1962_4406.t58 VSS 0.02309f
C529 a_n1962_4406.n116 VSS 0.05185f
C530 a_n1962_4406.n117 VSS 0.20376f
C531 a_n1962_4406.t47 VSS 0.02309f
C532 a_n1962_4406.t99 VSS 0.02309f
C533 a_n1962_4406.n118 VSS 0.05185f
C534 a_n1962_4406.n119 VSS 0.20376f
C535 a_n1962_4406.n120 VSS 0.20376f
C536 a_n1962_4406.n121 VSS 0.05185f
C537 a_n1962_4406.t59 VSS 0.02309f
C538 VOUT.n0 VSS 0.0137f
C539 VOUT.n1 VSS 0.01337f
C540 VOUT.n2 VSS 0.11544f
C541 VOUT.n3 VSS 0.01337f
C542 VOUT.n4 VSS 0.05946f
C543 VOUT.n5 VSS 0.01337f
C544 VOUT.n6 VSS 0.05946f
C545 VOUT.n7 VSS 0.01337f
C546 VOUT.n8 VSS 0.05946f
C547 VOUT.n9 VSS 0.01337f
C548 VOUT.n10 VSS 0.05946f
C549 VOUT.n11 VSS 0.01337f
C550 VOUT.n12 VSS 0.06305f
C551 VOUT.n13 VSS 0.0137f
C552 VOUT.n14 VSS 0.01337f
C553 VOUT.n15 VSS 0.11544f
C554 VOUT.n16 VSS 0.01337f
C555 VOUT.n17 VSS 0.05946f
C556 VOUT.n18 VSS 0.01337f
C557 VOUT.n19 VSS 0.05946f
C558 VOUT.n20 VSS 0.01337f
C559 VOUT.n21 VSS 0.05946f
C560 VOUT.n22 VSS 0.01337f
C561 VOUT.n23 VSS 0.05946f
C562 VOUT.n24 VSS 0.01337f
C563 VOUT.n25 VSS 0.06305f
C564 VOUT.n26 VSS 0.01996f
C565 VOUT.n27 VSS 0.01873f
C566 VOUT.n28 VSS 0.42323f
C567 VOUT.n29 VSS 0.01873f
C568 VOUT.n30 VSS 0.21781f
C569 VOUT.n31 VSS 0.02082f
C570 VOUT.n32 VSS 0.01873f
C571 VOUT.n33 VSS 0.46347f
C572 VOUT.n34 VSS 0.01873f
C573 VOUT.n35 VSS 0.21781f
C574 VOUT.n36 VSS 0.02009f
C575 VOUT.n37 VSS 0.01873f
C576 VOUT.n38 VSS 0.38202f
C577 VOUT.n39 VSS 0.01873f
C578 VOUT.n40 VSS 0.25889f
C579 VOUT.n41 VSS 0.02082f
C580 VOUT.n42 VSS 0.01873f
C581 VOUT.n43 VSS 0.46347f
C582 VOUT.n44 VSS 0.01873f
C583 VOUT.n45 VSS 0.21781f
C584 VOUT.n46 VSS 0.02009f
C585 VOUT.n47 VSS 0.01873f
C586 VOUT.n48 VSS 0.38202f
C587 VOUT.n49 VSS 0.01873f
C588 VOUT.n50 VSS 0.25889f
C589 VOUT.n51 VSS 0.02082f
C590 VOUT.n52 VSS 0.01873f
C591 VOUT.n53 VSS 0.46347f
C592 VOUT.n54 VSS 0.01873f
C593 VOUT.n55 VSS 0.21781f
C594 VOUT.n56 VSS 0.02009f
C595 VOUT.n57 VSS 0.01873f
C596 VOUT.n58 VSS 0.38202f
C597 VOUT.n59 VSS 0.01873f
C598 VOUT.n60 VSS 0.25889f
C599 VOUT.n61 VSS 0.02082f
C600 VOUT.n62 VSS 0.01873f
C601 VOUT.n63 VSS 0.46347f
C602 VOUT.n64 VSS 0.01873f
C603 VOUT.n65 VSS 0.21781f
C604 VOUT.n66 VSS 0.02009f
C605 VOUT.n67 VSS 0.01873f
C606 VOUT.n68 VSS 0.38202f
C607 VOUT.n69 VSS 0.01873f
C608 VOUT.n70 VSS 0.25889f
C609 VOUT.n71 VSS 0.01923f
C610 VOUT.n72 VSS 0.01873f
C611 VOUT.n73 VSS 0.25961f
C612 VOUT.n74 VSS 0.01873f
C613 VOUT.n75 VSS 0.29916f
C614 VOUT.n76 VSS 0.3698f
C615 VOUT.n77 VSS 0.13857f
C616 VOUT.n78 VSS 0.17966f
C617 VOUT.n79 VSS 0.13857f
C618 VOUT.n80 VSS 0.17966f
C619 VOUT.n81 VSS 0.13857f
C620 VOUT.n82 VSS 0.17966f
C621 VOUT.n83 VSS 0.13857f
C622 VOUT.n84 VSS 0.28975f
C623 VOUT.t78 VSS 0.17711p
C624 VOUT.n85 VSS 59.9272f
C625 VOUT.n86 VSS 0.4653f
C626 VOUT.n87 VSS 0.3048f
C627 a_3868_4185.t0 VSS 0.01921f
C628 a_3868_4185.t17 VSS 0.01921f
C629 a_3868_4185.t16 VSS 0.01921f
C630 a_3868_4185.n0 VSS 0.04532f
C631 a_3868_4185.t28 VSS 0.01921f
C632 a_3868_4185.t73 VSS 0.01921f
C633 a_3868_4185.n1 VSS 0.04313f
C634 a_3868_4185.n2 VSS 0.30359f
C635 a_3868_4185.t62 VSS 0.01921f
C636 a_3868_4185.t5 VSS 0.01921f
C637 a_3868_4185.n3 VSS 0.04313f
C638 a_3868_4185.n4 VSS 0.16949f
C639 a_3868_4185.t27 VSS 0.01921f
C640 a_3868_4185.t70 VSS 0.01921f
C641 a_3868_4185.n5 VSS 0.04313f
C642 a_3868_4185.n6 VSS 0.16949f
C643 a_3868_4185.t61 VSS 0.01921f
C644 a_3868_4185.t4 VSS 0.01921f
C645 a_3868_4185.n7 VSS 0.04313f
C646 a_3868_4185.n8 VSS 0.16949f
C647 a_3868_4185.t11 VSS 0.01921f
C648 a_3868_4185.t65 VSS 0.01921f
C649 a_3868_4185.n9 VSS 0.04313f
C650 a_3868_4185.n10 VSS 0.16949f
C651 a_3868_4185.t79 VSS 0.01921f
C652 a_3868_4185.t31 VSS 0.01921f
C653 a_3868_4185.n11 VSS 0.04313f
C654 a_3868_4185.n12 VSS 0.16949f
C655 a_3868_4185.t33 VSS 0.01921f
C656 a_3868_4185.t1 VSS 0.01921f
C657 a_3868_4185.n13 VSS 0.04532f
C658 a_3868_4185.t59 VSS 0.01921f
C659 a_3868_4185.t15 VSS 0.01921f
C660 a_3868_4185.n14 VSS 0.04313f
C661 a_3868_4185.n15 VSS 0.30359f
C662 a_3868_4185.t22 VSS 0.01921f
C663 a_3868_4185.t78 VSS 0.01921f
C664 a_3868_4185.n16 VSS 0.04313f
C665 a_3868_4185.n17 VSS 0.16949f
C666 a_3868_4185.t58 VSS 0.01921f
C667 a_3868_4185.t14 VSS 0.01921f
C668 a_3868_4185.n18 VSS 0.04313f
C669 a_3868_4185.n19 VSS 0.16949f
C670 a_3868_4185.t21 VSS 0.01921f
C671 a_3868_4185.t77 VSS 0.01921f
C672 a_3868_4185.n20 VSS 0.04313f
C673 a_3868_4185.n21 VSS 0.16949f
C674 a_3868_4185.t74 VSS 0.01921f
C675 a_3868_4185.t36 VSS 0.01921f
C676 a_3868_4185.n22 VSS 0.04313f
C677 a_3868_4185.n23 VSS 0.16949f
C678 a_3868_4185.t9 VSS 0.01921f
C679 a_3868_4185.t67 VSS 0.01921f
C680 a_3868_4185.n24 VSS 0.04313f
C681 a_3868_4185.n25 VSS 0.16949f
C682 a_3868_4185.t18 VSS 0.01921f
C683 a_3868_4185.t29 VSS 0.01921f
C684 a_3868_4185.n26 VSS 0.04313f
C685 a_3868_4185.n27 VSS 0.15383f
C686 a_3868_4185.t51 VSS 0.01921f
C687 a_3868_4185.t34 VSS 0.01921f
C688 a_3868_4185.n28 VSS 0.04532f
C689 a_3868_4185.t55 VSS 0.01921f
C690 a_3868_4185.t63 VSS 0.01921f
C691 a_3868_4185.n29 VSS 0.04313f
C692 a_3868_4185.n30 VSS 0.30359f
C693 a_3868_4185.t46 VSS 0.01921f
C694 a_3868_4185.t25 VSS 0.01921f
C695 a_3868_4185.n31 VSS 0.04313f
C696 a_3868_4185.n32 VSS 0.16949f
C697 a_3868_4185.t54 VSS 0.01921f
C698 a_3868_4185.t60 VSS 0.01921f
C699 a_3868_4185.n33 VSS 0.04313f
C700 a_3868_4185.n34 VSS 0.16949f
C701 a_3868_4185.t45 VSS 0.01921f
C702 a_3868_4185.t26 VSS 0.01921f
C703 a_3868_4185.n35 VSS 0.04313f
C704 a_3868_4185.n36 VSS 0.16949f
C705 a_3868_4185.t48 VSS 0.01921f
C706 a_3868_4185.t76 VSS 0.01921f
C707 a_3868_4185.n37 VSS 0.04313f
C708 a_3868_4185.n38 VSS 0.16949f
C709 a_3868_4185.t40 VSS 0.01921f
C710 a_3868_4185.t10 VSS 0.01921f
C711 a_3868_4185.n39 VSS 0.04313f
C712 a_3868_4185.n40 VSS 0.16949f
C713 a_3868_4185.t44 VSS 0.01921f
C714 a_3868_4185.t19 VSS 0.01921f
C715 a_3868_4185.n41 VSS 0.04313f
C716 a_3868_4185.n42 VSS 0.23792f
C717 a_3868_4185.n43 VSS 0.2626f
C718 a_3868_4185.t13 VSS 0.01921f
C719 a_3868_4185.t12 VSS 0.01921f
C720 a_3868_4185.n44 VSS 0.04532f
C721 a_3868_4185.t69 VSS 0.01921f
C722 a_3868_4185.t24 VSS 0.01921f
C723 a_3868_4185.n45 VSS 0.04313f
C724 a_3868_4185.n46 VSS 0.30359f
C725 a_3868_4185.t3 VSS 0.01921f
C726 a_3868_4185.t57 VSS 0.01921f
C727 a_3868_4185.n47 VSS 0.04313f
C728 a_3868_4185.n48 VSS 0.16949f
C729 a_3868_4185.t68 VSS 0.01921f
C730 a_3868_4185.t23 VSS 0.01921f
C731 a_3868_4185.n49 VSS 0.04313f
C732 a_3868_4185.n50 VSS 0.16949f
C733 a_3868_4185.t2 VSS 0.01921f
C734 a_3868_4185.t56 VSS 0.01921f
C735 a_3868_4185.n51 VSS 0.04313f
C736 a_3868_4185.n52 VSS 0.16949f
C737 a_3868_4185.t64 VSS 0.01921f
C738 a_3868_4185.t8 VSS 0.01921f
C739 a_3868_4185.n53 VSS 0.04313f
C740 a_3868_4185.n54 VSS 0.16949f
C741 a_3868_4185.t30 VSS 0.01921f
C742 a_3868_4185.t75 VSS 0.01921f
C743 a_3868_4185.n55 VSS 0.04313f
C744 a_3868_4185.n56 VSS 0.16949f
C745 a_3868_4185.t38 VSS 0.01921f
C746 a_3868_4185.t37 VSS 0.01921f
C747 a_3868_4185.n57 VSS 0.04313f
C748 a_3868_4185.n58 VSS 0.15383f
C749 a_3868_4185.t35 VSS 0.01921f
C750 a_3868_4185.t53 VSS 0.01921f
C751 a_3868_4185.n59 VSS 0.04532f
C752 a_3868_4185.t7 VSS 0.01921f
C753 a_3868_4185.t42 VSS 0.01921f
C754 a_3868_4185.n60 VSS 0.04313f
C755 a_3868_4185.n61 VSS 0.30359f
C756 a_3868_4185.t72 VSS 0.01921f
C757 a_3868_4185.t50 VSS 0.01921f
C758 a_3868_4185.n62 VSS 0.04313f
C759 a_3868_4185.n63 VSS 0.16949f
C760 a_3868_4185.t6 VSS 0.01921f
C761 a_3868_4185.t41 VSS 0.01921f
C762 a_3868_4185.n64 VSS 0.04313f
C763 a_3868_4185.n65 VSS 0.16949f
C764 a_3868_4185.t71 VSS 0.01921f
C765 a_3868_4185.t49 VSS 0.01921f
C766 a_3868_4185.n66 VSS 0.04313f
C767 a_3868_4185.n67 VSS 0.16949f
C768 a_3868_4185.t32 VSS 0.01921f
C769 a_3868_4185.t52 VSS 0.01921f
C770 a_3868_4185.n68 VSS 0.04313f
C771 a_3868_4185.n69 VSS 0.16949f
C772 a_3868_4185.t66 VSS 0.01921f
C773 a_3868_4185.t43 VSS 0.01921f
C774 a_3868_4185.n70 VSS 0.04313f
C775 a_3868_4185.n71 VSS 0.16949f
C776 a_3868_4185.t20 VSS 0.01921f
C777 a_3868_4185.t47 VSS 0.01921f
C778 a_3868_4185.n72 VSS 0.04313f
C779 a_3868_4185.n73 VSS 0.23792f
C780 a_3868_4185.n74 VSS 0.2626f
C781 a_3868_4185.n75 VSS 0.20915f
C782 a_3868_4185.n76 VSS 0.15383f
C783 a_3868_4185.n77 VSS 0.04313f
C784 a_3868_4185.t39 VSS 0.01921f
C785 a_3329_8823.t32 VSS 0.01153f
C786 a_3329_8823.t24 VSS 0.01153f
C787 a_3329_8823.t9 VSS 0.01153f
C788 a_3329_8823.n0 VSS 0.03611f
C789 a_3329_8823.t15 VSS 0.01153f
C790 a_3329_8823.t33 VSS 0.01153f
C791 a_3329_8823.n1 VSS 0.03366f
C792 a_3329_8823.n2 VSS 0.73879f
C793 a_3329_8823.t36 VSS 0.01153f
C794 a_3329_8823.t27 VSS 0.01153f
C795 a_3329_8823.n3 VSS 0.03741f
C796 a_3329_8823.t34 VSS 0.01153f
C797 a_3329_8823.t30 VSS 0.01153f
C798 a_3329_8823.n4 VSS 0.03366f
C799 a_3329_8823.n5 VSS 0.81133f
C800 a_3329_8823.t4 VSS 0.01153f
C801 a_3329_8823.t2 VSS 0.01153f
C802 a_3329_8823.n6 VSS 0.03456f
C803 a_3329_8823.t31 VSS 0.01153f
C804 a_3329_8823.t16 VSS 0.01153f
C805 a_3329_8823.n7 VSS 0.03366f
C806 a_3329_8823.n8 VSS 0.46658f
C807 a_3329_8823.t21 VSS 0.01153f
C808 a_3329_8823.t23 VSS 0.01153f
C809 a_3329_8823.n9 VSS 0.03366f
C810 a_3329_8823.n10 VSS 0.26536f
C811 a_3329_8823.t10 VSS 0.01153f
C812 a_3329_8823.t35 VSS 0.01153f
C813 a_3329_8823.n11 VSS 0.03366f
C814 a_3329_8823.n12 VSS 0.3176f
C815 a_3329_8823.t47 VSS 0.01153f
C816 a_3329_8823.t43 VSS 0.01153f
C817 a_3329_8823.n13 VSS 0.0272f
C818 a_3329_8823.t64 VSS 0.01153f
C819 a_3329_8823.t76 VSS 0.01153f
C820 a_3329_8823.n14 VSS 0.02589f
C821 a_3329_8823.n15 VSS 0.18219f
C822 a_3329_8823.t56 VSS 0.01153f
C823 a_3329_8823.t65 VSS 0.01153f
C824 a_3329_8823.n16 VSS 0.02589f
C825 a_3329_8823.n17 VSS 0.10172f
C826 a_3329_8823.t70 VSS 0.01153f
C827 a_3329_8823.t75 VSS 0.01153f
C828 a_3329_8823.n18 VSS 0.02589f
C829 a_3329_8823.n19 VSS 0.10208f
C830 a_3329_8823.t40 VSS 0.01153f
C831 a_3329_8823.t45 VSS 0.01153f
C832 a_3329_8823.n20 VSS 0.02589f
C833 a_3329_8823.n21 VSS 0.07415f
C834 a_3329_8823.t78 VSS 0.01153f
C835 a_3329_8823.t50 VSS 0.01153f
C836 a_3329_8823.n22 VSS 0.02742f
C837 a_3329_8823.t62 VSS 0.01153f
C838 a_3329_8823.t48 VSS 0.01153f
C839 a_3329_8823.n23 VSS 0.02589f
C840 a_3329_8823.n24 VSS 0.19587f
C841 a_3329_8823.t69 VSS 0.01153f
C842 a_3329_8823.t53 VSS 0.01153f
C843 a_3329_8823.n25 VSS 0.02589f
C844 a_3329_8823.n26 VSS 0.10208f
C845 a_3329_8823.t57 VSS 0.01153f
C846 a_3329_8823.t52 VSS 0.01153f
C847 a_3329_8823.n27 VSS 0.02589f
C848 a_3329_8823.n28 VSS 0.12674f
C849 a_3329_8823.n29 VSS 0.10458f
C850 a_3329_8823.t72 VSS 0.01153f
C851 a_3329_8823.t60 VSS 0.01153f
C852 a_3329_8823.n30 VSS 0.02589f
C853 a_3329_8823.n31 VSS 0.09175f
C854 a_3329_8823.t68 VSS 0.01153f
C855 a_3329_8823.t77 VSS 0.01153f
C856 a_3329_8823.n32 VSS 0.0272f
C857 a_3329_8823.t74 VSS 0.01153f
C858 a_3329_8823.t66 VSS 0.01153f
C859 a_3329_8823.n33 VSS 0.02589f
C860 a_3329_8823.n34 VSS 0.18219f
C861 a_3329_8823.t46 VSS 0.01153f
C862 a_3329_8823.t59 VSS 0.01153f
C863 a_3329_8823.n35 VSS 0.02589f
C864 a_3329_8823.n36 VSS 0.10172f
C865 a_3329_8823.t41 VSS 0.01153f
C866 a_3329_8823.t42 VSS 0.01153f
C867 a_3329_8823.n37 VSS 0.02589f
C868 a_3329_8823.n38 VSS 0.10208f
C869 a_3329_8823.t44 VSS 0.01153f
C870 a_3329_8823.t61 VSS 0.01153f
C871 a_3329_8823.n39 VSS 0.02589f
C872 a_3329_8823.n40 VSS 0.07415f
C873 a_3329_8823.t49 VSS 0.01153f
C874 a_3329_8823.t58 VSS 0.01153f
C875 a_3329_8823.n41 VSS 0.02746f
C876 a_3329_8823.t51 VSS 0.01153f
C877 a_3329_8823.t79 VSS 0.01153f
C878 a_3329_8823.n42 VSS 0.02589f
C879 a_3329_8823.n43 VSS 0.1982f
C880 a_3329_8823.t55 VSS 0.01153f
C881 a_3329_8823.t63 VSS 0.01153f
C882 a_3329_8823.n44 VSS 0.02589f
C883 a_3329_8823.n45 VSS 0.10208f
C884 a_3329_8823.t54 VSS 0.01153f
C885 a_3329_8823.t71 VSS 0.01153f
C886 a_3329_8823.n46 VSS 0.02589f
C887 a_3329_8823.n47 VSS 0.12674f
C888 a_3329_8823.n48 VSS 0.10458f
C889 a_3329_8823.t73 VSS 0.01153f
C890 a_3329_8823.t67 VSS 0.01153f
C891 a_3329_8823.n49 VSS 0.02589f
C892 a_3329_8823.n50 VSS 0.21634f
C893 a_3329_8823.n51 VSS 0.38602f
C894 a_3329_8823.n52 VSS 0.42211f
C895 a_3329_8823.n53 VSS 0.24874f
C896 a_3329_8823.n54 VSS 0.32288f
C897 a_3329_8823.t14 VSS 0.01153f
C898 a_3329_8823.t13 VSS 0.01153f
C899 a_3329_8823.n55 VSS 0.03611f
C900 a_3329_8823.t37 VSS 0.01153f
C901 a_3329_8823.t20 VSS 0.01153f
C902 a_3329_8823.n56 VSS 0.03366f
C903 a_3329_8823.n57 VSS 0.73879f
C904 a_3329_8823.t17 VSS 0.01153f
C905 a_3329_8823.t7 VSS 0.01153f
C906 a_3329_8823.n58 VSS 0.03741f
C907 a_3329_8823.t26 VSS 0.01153f
C908 a_3329_8823.t28 VSS 0.01153f
C909 a_3329_8823.n59 VSS 0.03366f
C910 a_3329_8823.n60 VSS 0.81133f
C911 a_3329_8823.t3 VSS 0.01153f
C912 a_3329_8823.t29 VSS 0.01153f
C913 a_3329_8823.n61 VSS 0.03611f
C914 a_3329_8823.t11 VSS 0.01153f
C915 a_3329_8823.t12 VSS 0.01153f
C916 a_3329_8823.n62 VSS 0.03366f
C917 a_3329_8823.n63 VSS 0.73879f
C918 a_3329_8823.t25 VSS 0.01153f
C919 a_3329_8823.t6 VSS 0.01153f
C920 a_3329_8823.n64 VSS 0.03456f
C921 a_3329_8823.t18 VSS 0.01153f
C922 a_3329_8823.t19 VSS 0.01153f
C923 a_3329_8823.n65 VSS 0.03366f
C924 a_3329_8823.n66 VSS 0.46658f
C925 a_3329_8823.t39 VSS 0.01153f
C926 a_3329_8823.t38 VSS 0.01153f
C927 a_3329_8823.n67 VSS 0.03366f
C928 a_3329_8823.n68 VSS 0.26536f
C929 a_3329_8823.t8 VSS 0.01153f
C930 a_3329_8823.t1 VSS 0.01153f
C931 a_3329_8823.n69 VSS 0.03366f
C932 a_3329_8823.n70 VSS 0.38027f
C933 a_3329_8823.n71 VSS 0.45864f
C934 a_3329_8823.n72 VSS 0.24903f
C935 a_3329_8823.n73 VSS 0.32288f
C936 a_3329_8823.n74 VSS 0.24903f
C937 a_3329_8823.t5 VSS 0.01153f
C938 a_3329_8823.t22 VSS 0.01153f
C939 a_3329_8823.n75 VSS 0.03366f
C940 a_3329_8823.n76 VSS 0.81133f
C941 a_3329_8823.n77 VSS 0.03741f
C942 a_3329_8823.t0 VSS 0.01153f
C943 IBIAS.t5 VSS 0.02161f
C944 IBIAS.t8 VSS 0.02161f
C945 IBIAS.n0 VSS 0.05408f
C946 IBIAS.t4 VSS 0.25108f
C947 IBIAS.n1 VSS 0.51806f
C948 IBIAS.t6 VSS 0.25108f
C949 IBIAS.n2 VSS 0.22293f
C950 IBIAS.t1 VSS 0.02161f
C951 IBIAS.t7 VSS 0.02161f
C952 IBIAS.n3 VSS 0.05318f
C953 IBIAS.n4 VSS 0.31686f
C954 IBIAS.t0 VSS 0.25108f
C955 IBIAS.n5 VSS 0.22293f
C956 IBIAS.t2 VSS 0.25108f
C957 IBIAS.n6 VSS 0.22293f
C958 IBIAS.t9 VSS 0.02161f
C959 IBIAS.t3 VSS 0.02161f
C960 IBIAS.n7 VSS 0.05318f
C961 IBIAS.n8 VSS 0.41073f
C962 IBIAS.t42 VSS 0.2525f
C963 IBIAS.t69 VSS 0.25121f
C964 IBIAS.n9 VSS 0.50883f
C965 IBIAS.t102 VSS 0.25121f
C966 IBIAS.n10 VSS 0.26494f
C967 IBIAS.t19 VSS 0.25121f
C968 IBIAS.n11 VSS 0.26494f
C969 IBIAS.t16 VSS 0.25121f
C970 IBIAS.n12 VSS 0.26494f
C971 IBIAS.t38 VSS 0.25121f
C972 IBIAS.n13 VSS 0.69526f
C973 IBIAS.t20 VSS 0.2525f
C974 IBIAS.t21 VSS 0.25121f
C975 IBIAS.n14 VSS 0.60881f
C976 IBIAS.t58 VSS 0.25121f
C977 IBIAS.n15 VSS 0.36492f
C978 IBIAS.t66 VSS 0.25121f
C979 IBIAS.n16 VSS 0.36492f
C980 IBIAS.t64 VSS 0.25121f
C981 IBIAS.n17 VSS 0.36492f
C982 IBIAS.t89 VSS 0.25121f
C983 IBIAS.n18 VSS 0.5303f
C984 IBIAS.n19 VSS 0.84775f
C985 IBIAS.t46 VSS 0.25355f
C986 IBIAS.t72 VSS 0.25121f
C987 IBIAS.n20 VSS 0.80771f
C988 IBIAS.t17 VSS 0.25121f
C989 IBIAS.n21 VSS 0.36492f
C990 IBIAS.t39 VSS 0.25121f
C991 IBIAS.n22 VSS 0.36492f
C992 IBIAS.t37 VSS 0.25121f
C993 IBIAS.n23 VSS 0.36492f
C994 IBIAS.t35 VSS 0.25121f
C995 IBIAS.n24 VSS 0.43024f
C996 IBIAS.n25 VSS 0.36752f
C997 IBIAS.t40 VSS 0.2525f
C998 IBIAS.t43 VSS 0.25121f
C999 IBIAS.n26 VSS 0.60881f
C1000 IBIAS.t83 VSS 0.25121f
C1001 IBIAS.n27 VSS 0.36492f
C1002 IBIAS.t91 VSS 0.25121f
C1003 IBIAS.n28 VSS 0.36492f
C1004 IBIAS.t90 VSS 0.25121f
C1005 IBIAS.n29 VSS 0.36492f
C1006 IBIAS.t18 VSS 0.25121f
C1007 IBIAS.n30 VSS 0.5303f
C1008 IBIAS.n31 VSS 0.46741f
C1009 IBIAS.t74 VSS 0.25355f
C1010 IBIAS.t104 VSS 0.25121f
C1011 IBIAS.n32 VSS 0.80771f
C1012 IBIAS.t44 VSS 0.25121f
C1013 IBIAS.n33 VSS 0.36492f
C1014 IBIAS.t65 VSS 0.25121f
C1015 IBIAS.n34 VSS 0.36492f
C1016 IBIAS.t63 VSS 0.25121f
C1017 IBIAS.n35 VSS 0.36492f
C1018 IBIAS.t62 VSS 0.25121f
C1019 IBIAS.n36 VSS 0.43024f
C1020 IBIAS.n37 VSS 0.36752f
C1021 IBIAS.t70 VSS 0.2525f
C1022 IBIAS.t75 VSS 0.25121f
C1023 IBIAS.n38 VSS 0.60881f
C1024 IBIAS.t11 VSS 0.25121f
C1025 IBIAS.n39 VSS 0.36492f
C1026 IBIAS.t25 VSS 0.25121f
C1027 IBIAS.n40 VSS 0.36492f
C1028 IBIAS.t22 VSS 0.25121f
C1029 IBIAS.n41 VSS 0.36492f
C1030 IBIAS.t47 VSS 0.25121f
C1031 IBIAS.n42 VSS 0.5303f
C1032 IBIAS.n43 VSS 0.46741f
C1033 IBIAS.t108 VSS 0.25355f
C1034 IBIAS.t32 VSS 0.25121f
C1035 IBIAS.n44 VSS 0.80771f
C1036 IBIAS.t76 VSS 0.25121f
C1037 IBIAS.n45 VSS 0.36492f
C1038 IBIAS.t98 VSS 0.25121f
C1039 IBIAS.n46 VSS 0.36492f
C1040 IBIAS.t96 VSS 0.25121f
C1041 IBIAS.n47 VSS 0.36492f
C1042 IBIAS.t93 VSS 0.25121f
C1043 IBIAS.n48 VSS 0.43024f
C1044 IBIAS.n49 VSS 0.36752f
C1045 IBIAS.t73 VSS 0.2525f
C1046 IBIAS.t79 VSS 0.25121f
C1047 IBIAS.n50 VSS 0.60881f
C1048 IBIAS.t12 VSS 0.25121f
C1049 IBIAS.n51 VSS 0.36492f
C1050 IBIAS.t26 VSS 0.25121f
C1051 IBIAS.n52 VSS 0.36492f
C1052 IBIAS.t24 VSS 0.25121f
C1053 IBIAS.n53 VSS 0.36492f
C1054 IBIAS.t48 VSS 0.25121f
C1055 IBIAS.n54 VSS 0.5303f
C1056 IBIAS.n55 VSS 0.46741f
C1057 IBIAS.t109 VSS 0.25355f
C1058 IBIAS.t33 VSS 0.25121f
C1059 IBIAS.n56 VSS 0.80771f
C1060 IBIAS.t77 VSS 0.25121f
C1061 IBIAS.n57 VSS 0.36492f
C1062 IBIAS.t99 VSS 0.25121f
C1063 IBIAS.n58 VSS 0.36492f
C1064 IBIAS.t97 VSS 0.25121f
C1065 IBIAS.n59 VSS 0.36492f
C1066 IBIAS.t94 VSS 0.25121f
C1067 IBIAS.n60 VSS 0.43024f
C1068 IBIAS.n61 VSS 0.36752f
C1069 IBIAS.t34 VSS 0.25461f
C1070 IBIAS.t51 VSS 0.25121f
C1071 IBIAS.n62 VSS 0.90663f
C1072 IBIAS.t49 VSS 0.25121f
C1073 IBIAS.n63 VSS 0.26494f
C1074 IBIAS.t67 VSS 0.25121f
C1075 IBIAS.n64 VSS 0.26494f
C1076 IBIAS.t50 VSS 0.25121f
C1077 IBIAS.n65 VSS 0.26494f
C1078 IBIAS.t68 VSS 0.25121f
C1079 IBIAS.n66 VSS 0.5303f
C1080 IBIAS.n67 VSS 1.63924f
C1081 IBIAS.t60 VSS 0.2525f
C1082 IBIAS.t61 VSS 0.25121f
C1083 IBIAS.n68 VSS 0.50883f
C1084 IBIAS.t36 VSS 0.25121f
C1085 IBIAS.n69 VSS 0.26494f
C1086 IBIAS.t107 VSS 0.25121f
C1087 IBIAS.n70 VSS 0.26494f
C1088 IBIAS.t10 VSS 0.25121f
C1089 IBIAS.n71 VSS 0.26494f
C1090 IBIAS.t13 VSS 0.25121f
C1091 IBIAS.n72 VSS 0.26494f
C1092 IBIAS.t14 VSS 0.25121f
C1093 IBIAS.n73 VSS 0.26494f
C1094 IBIAS.t59 VSS 0.25121f
C1095 IBIAS.n74 VSS 0.42805f
C1096 IBIAS.t86 VSS 0.2525f
C1097 IBIAS.t87 VSS 0.25121f
C1098 IBIAS.n75 VSS 0.60881f
C1099 IBIAS.t30 VSS 0.25121f
C1100 IBIAS.n76 VSS 0.36492f
C1101 IBIAS.t31 VSS 0.25121f
C1102 IBIAS.n77 VSS 0.528f
C1103 IBIAS.t15 VSS 0.25355f
C1104 IBIAS.t85 VSS 0.25121f
C1105 IBIAS.n78 VSS 0.80771f
C1106 IBIAS.t88 VSS 0.25121f
C1107 IBIAS.n79 VSS 0.36492f
C1108 IBIAS.t29 VSS 0.25121f
C1109 IBIAS.n80 VSS 0.42798f
C1110 IBIAS.t52 VSS 0.2525f
C1111 IBIAS.t57 VSS 0.25121f
C1112 IBIAS.n81 VSS 0.60881f
C1113 IBIAS.t101 VSS 0.25121f
C1114 IBIAS.n82 VSS 0.36492f
C1115 IBIAS.t105 VSS 0.25121f
C1116 IBIAS.n83 VSS 0.528f
C1117 IBIAS.t81 VSS 0.25355f
C1118 IBIAS.t45 VSS 0.25121f
C1119 IBIAS.n84 VSS 0.80771f
C1120 IBIAS.t55 VSS 0.25121f
C1121 IBIAS.n85 VSS 0.36492f
C1122 IBIAS.t95 VSS 0.25121f
C1123 IBIAS.n86 VSS 0.42798f
C1124 IBIAS.t53 VSS 0.2525f
C1125 IBIAS.t56 VSS 0.25121f
C1126 IBIAS.n87 VSS 0.60881f
C1127 IBIAS.t100 VSS 0.25121f
C1128 IBIAS.n88 VSS 0.36492f
C1129 IBIAS.t103 VSS 0.25121f
C1130 IBIAS.n89 VSS 0.528f
C1131 IBIAS.t80 VSS 0.25355f
C1132 IBIAS.t41 VSS 0.25121f
C1133 IBIAS.n90 VSS 0.80771f
C1134 IBIAS.t54 VSS 0.25121f
C1135 IBIAS.n91 VSS 0.36492f
C1136 IBIAS.t92 VSS 0.25121f
C1137 IBIAS.n92 VSS 0.42798f
C1138 IBIAS.t27 VSS 0.2525f
C1139 IBIAS.t28 VSS 0.25134f
C1140 IBIAS.n93 VSS 0.51568f
C1141 IBIAS.t106 VSS 0.25134f
C1142 IBIAS.n94 VSS 0.27179f
C1143 IBIAS.t71 VSS 0.25134f
C1144 IBIAS.n95 VSS 0.27179f
C1145 IBIAS.t78 VSS 0.25134f
C1146 IBIAS.n96 VSS 0.27179f
C1147 IBIAS.t82 VSS 0.25134f
C1148 IBIAS.n97 VSS 0.27179f
C1149 IBIAS.t84 VSS 0.25134f
C1150 IBIAS.n98 VSS 0.27179f
C1151 IBIAS.t23 VSS 0.25121f
C1152 IBIAS.n99 VSS 0.51945f
C1153 IBIAS.n100 VSS 0.6264f
C1154 IBIAS.n101 VSS 0.46851f
C1155 IBIAS.n102 VSS 0.36859f
C1156 IBIAS.n103 VSS 0.46851f
C1157 IBIAS.n104 VSS 0.36859f
C1158 IBIAS.n105 VSS 0.46858f
C1159 IBIAS.n106 VSS 0.44083f
C1160 IBIAS.n107 VSS 3.49898f
C1161 IBIAS.n108 VSS 2.57679f
C1162 VDD.n0 VSS 0.02345f
C1163 VDD.n1 VSS 0.01701f
C1164 VDD.t79 VSS 0.01949f
C1165 VDD.n3 VSS 0.01858f
C1166 VDD.n4 VSS 0.0147f
C1167 VDD.n5 VSS 0.01701f
C1168 VDD.n6 VSS 0.0147f
C1169 VDD.t72 VSS 0.01949f
C1170 VDD.n8 VSS 0.01858f
C1171 VDD.n9 VSS 0.0147f
C1172 VDD.n10 VSS 0.01701f
C1173 VDD.n11 VSS 0.0147f
C1174 VDD.t90 VSS 0.01949f
C1175 VDD.n13 VSS 0.01858f
C1176 VDD.n14 VSS 0.0147f
C1177 VDD.n15 VSS 0.01701f
C1178 VDD.n16 VSS 0.0147f
C1179 VDD.t77 VSS 0.01949f
C1180 VDD.n18 VSS 0.01858f
C1181 VDD.n19 VSS 0.0147f
C1182 VDD.n20 VSS 0.01701f
C1183 VDD.n21 VSS 0.0147f
C1184 VDD.t83 VSS 0.01949f
C1185 VDD.n23 VSS 0.01858f
C1186 VDD.n24 VSS 0.0147f
C1187 VDD.n25 VSS 0.01701f
C1188 VDD.n26 VSS 0.0147f
C1189 VDD.t92 VSS 0.01949f
C1190 VDD.n28 VSS 0.01858f
C1191 VDD.n29 VSS 0.0147f
C1192 VDD.n30 VSS 0.02306f
C1193 VDD.n31 VSS 0.0147f
C1194 VDD.t81 VSS 0.01949f
C1195 VDD.n33 VSS 0.02464f
C1196 VDD.n34 VSS 0.03911f
C1197 VDD.t80 VSS 0.09216f
C1198 VDD.n35 VSS 0.02588f
C1199 VDD.n36 VSS 0.0147f
C1200 VDD.n37 VSS 0.0147f
C1201 VDD.n38 VSS 0.02588f
C1202 VDD.t91 VSS 0.09216f
C1203 VDD.n39 VSS 0.02588f
C1204 VDD.n40 VSS 0.0147f
C1205 VDD.n41 VSS 0.0147f
C1206 VDD.n42 VSS 0.02588f
C1207 VDD.t82 VSS 0.09216f
C1208 VDD.n43 VSS 0.02588f
C1209 VDD.n44 VSS 0.0147f
C1210 VDD.n45 VSS 0.0147f
C1211 VDD.n46 VSS 0.02588f
C1212 VDD.t76 VSS 0.09216f
C1213 VDD.n47 VSS 0.02588f
C1214 VDD.n48 VSS 0.0147f
C1215 VDD.n49 VSS 0.0147f
C1216 VDD.n50 VSS 0.02588f
C1217 VDD.t89 VSS 0.09216f
C1218 VDD.n51 VSS 0.02588f
C1219 VDD.n52 VSS 0.0147f
C1220 VDD.n53 VSS 0.0147f
C1221 VDD.n54 VSS 0.02588f
C1222 VDD.t70 VSS 0.09216f
C1223 VDD.n55 VSS 0.02588f
C1224 VDD.n56 VSS 0.0147f
C1225 VDD.n57 VSS 0.0147f
C1226 VDD.n58 VSS 0.02588f
C1227 VDD.t78 VSS 0.09216f
C1228 VDD.n59 VSS 0.02588f
C1229 VDD.n60 VSS 0.01526f
C1230 VDD.n65 VSS 0.3162f
C1231 VDD.n69 VSS 0.3162f
C1232 VDD.n76 VSS 0.3162f
C1233 VDD.n83 VSS 0.3162f
C1234 VDD.n90 VSS 0.3162f
C1235 VDD.n97 VSS 0.52546f
C1236 VDD.t71 VSS 0.1581f
C1237 VDD.n126 VSS 0.37201f
C1238 VDD.n235 VSS 0.46036f
C1239 VDD.n243 VSS 0.19298f
C1240 VDD.n244 VSS 0.3162f
C1241 VDD.n250 VSS 0.28133f
C1242 VDD.n365 VSS 0.43711f
C1243 VDD.n366 VSS 0.28598f
C1244 VDD.t40 VSS 0.1581f
C1245 VDD.n367 VSS 0.18833f
C1246 VDD.n373 VSS 0.3162f
C1247 VDD.n374 VSS 0.25343f
C1248 VDD.t2 VSS 0.1581f
C1249 VDD.n375 VSS 0.22088f
C1250 VDD.n381 VSS 0.3162f
C1251 VDD.n382 VSS 0.22088f
C1252 VDD.t5 VSS 0.1581f
C1253 VDD.n383 VSS 0.25343f
C1254 VDD.n389 VSS 0.3162f
C1255 VDD.n390 VSS 0.18833f
C1256 VDD.t13 VSS 0.1581f
C1257 VDD.n391 VSS 0.28598f
C1258 VDD.n397 VSS 0.31388f
C1259 VDD.t15 VSS 0.1581f
C1260 VDD.n398 VSS 0.16043f
C1261 VDD.n399 VSS 0.3162f
C1262 VDD.n403 VSS 0.01078f
C1263 VDD.n406 VSS 0.07459f
C1264 VDD.n408 VSS 0.03842f
C1265 VDD.n410 VSS 0.03842f
C1266 VDD.n412 VSS 0.03842f
C1267 VDD.n414 VSS 0.03842f
C1268 VDD.n416 VSS 0.04074f
C1269 VDD.n417 VSS 0.02345f
C1270 VDD.t75 VSS 0.01535f
C1271 VDD.n418 VSS 0.01858f
C1272 VDD.n420 VSS 0.01701f
C1273 VDD.n421 VSS 0.0147f
C1274 VDD.t66 VSS 0.01535f
C1275 VDD.n422 VSS 0.01858f
C1276 VDD.n423 VSS 0.0147f
C1277 VDD.n425 VSS 0.01701f
C1278 VDD.n426 VSS 0.0147f
C1279 VDD.t63 VSS 0.01535f
C1280 VDD.n427 VSS 0.01858f
C1281 VDD.n428 VSS 0.0147f
C1282 VDD.n430 VSS 0.01701f
C1283 VDD.n431 VSS 0.0147f
C1284 VDD.t42 VSS 0.01535f
C1285 VDD.n432 VSS 0.01858f
C1286 VDD.n433 VSS 0.0147f
C1287 VDD.n435 VSS 0.01701f
C1288 VDD.n436 VSS 0.0147f
C1289 VDD.t57 VSS 0.01535f
C1290 VDD.n437 VSS 0.01858f
C1291 VDD.n438 VSS 0.0147f
C1292 VDD.n440 VSS 0.01701f
C1293 VDD.n441 VSS 0.0147f
C1294 VDD.t69 VSS 0.01535f
C1295 VDD.n442 VSS 0.01858f
C1296 VDD.n443 VSS 0.0147f
C1297 VDD.n445 VSS 0.01701f
C1298 VDD.n446 VSS 0.0147f
C1299 VDD.t52 VSS 0.01535f
C1300 VDD.n447 VSS 0.02464f
C1301 VDD.n448 VSS 0.0147f
C1302 VDD.n450 VSS 0.02306f
C1303 VDD.n451 VSS 0.03911f
C1304 VDD.t50 VSS 0.09216f
C1305 VDD.n452 VSS 0.02588f
C1306 VDD.n453 VSS 0.0147f
C1307 VDD.n454 VSS 0.0147f
C1308 VDD.n455 VSS 0.02588f
C1309 VDD.t67 VSS 0.09216f
C1310 VDD.n456 VSS 0.02588f
C1311 VDD.n457 VSS 0.0147f
C1312 VDD.n458 VSS 0.0147f
C1313 VDD.n459 VSS 0.02588f
C1314 VDD.t55 VSS 0.09216f
C1315 VDD.n460 VSS 0.02588f
C1316 VDD.n461 VSS 0.0147f
C1317 VDD.n462 VSS 0.0147f
C1318 VDD.n463 VSS 0.02588f
C1319 VDD.t39 VSS 0.09216f
C1320 VDD.n464 VSS 0.02588f
C1321 VDD.n465 VSS 0.0147f
C1322 VDD.n466 VSS 0.0147f
C1323 VDD.n467 VSS 0.02588f
C1324 VDD.t61 VSS 0.09216f
C1325 VDD.n468 VSS 0.02588f
C1326 VDD.n469 VSS 0.0147f
C1327 VDD.n470 VSS 0.0147f
C1328 VDD.n471 VSS 0.02588f
C1329 VDD.t64 VSS 0.09216f
C1330 VDD.n472 VSS 0.02588f
C1331 VDD.n473 VSS 0.0147f
C1332 VDD.n474 VSS 0.0147f
C1333 VDD.n475 VSS 0.02588f
C1334 VDD.t73 VSS 0.09216f
C1335 VDD.n476 VSS 0.02588f
C1336 VDD.n477 VSS 0.02345f
C1337 VDD.n480 VSS 0.07524f
C1338 VDD.n482 VSS 0.03842f
C1339 VDD.n484 VSS 0.0391f
C1340 VDD.n485 VSS 0.02184f
C1341 VDD.n486 VSS 0.01858f
C1342 VDD.n487 VSS 0.0147f
C1343 VDD.n488 VSS 0.01701f
C1344 VDD.n489 VSS 0.0147f
C1345 VDD.t45 VSS 0.01949f
C1346 VDD.n491 VSS 0.01858f
C1347 VDD.n492 VSS 0.0147f
C1348 VDD.n493 VSS 0.01701f
C1349 VDD.n494 VSS 0.0147f
C1350 VDD.t54 VSS 0.01949f
C1351 VDD.n496 VSS 0.01858f
C1352 VDD.n497 VSS 0.0147f
C1353 VDD.n498 VSS 0.02306f
C1354 VDD.n499 VSS 0.0147f
C1355 VDD.t88 VSS 0.01949f
C1356 VDD.n501 VSS 0.02464f
C1357 VDD.n502 VSS 0.03911f
C1358 VDD.t87 VSS 0.09216f
C1359 VDD.n503 VSS 0.02588f
C1360 VDD.n504 VSS 0.0147f
C1361 VDD.n505 VSS 0.0147f
C1362 VDD.n506 VSS 0.02588f
C1363 VDD.t53 VSS 0.09216f
C1364 VDD.n507 VSS 0.02588f
C1365 VDD.n508 VSS 0.0147f
C1366 VDD.n509 VSS 0.0147f
C1367 VDD.n510 VSS 0.02588f
C1368 VDD.t43 VSS 0.09216f
C1369 VDD.n511 VSS 0.02588f
C1370 VDD.n512 VSS 0.0147f
C1371 VDD.t97 VSS 0.01949f
C1372 VDD.n514 VSS 0.01701f
C1373 VDD.n515 VSS 0.0147f
C1374 VDD.n516 VSS 0.02588f
C1375 VDD.t96 VSS 0.09216f
C1376 VDD.n517 VSS 0.02588f
C1377 VDD.n518 VSS 0.04421f
C1378 VDD.n519 VSS 0.05881f
C1379 VDD.n520 VSS 0.04816f
C1380 VDD.n521 VSS 0.02184f
C1381 VDD.t86 VSS 0.01535f
C1382 VDD.n522 VSS 0.01858f
C1383 VDD.n524 VSS 0.01701f
C1384 VDD.n525 VSS 0.0147f
C1385 VDD.t49 VSS 0.01535f
C1386 VDD.n526 VSS 0.01858f
C1387 VDD.n527 VSS 0.0147f
C1388 VDD.n529 VSS 0.01701f
C1389 VDD.n530 VSS 0.0147f
C1390 VDD.t60 VSS 0.01535f
C1391 VDD.n531 VSS 0.01858f
C1392 VDD.n532 VSS 0.0147f
C1393 VDD.n534 VSS 0.01701f
C1394 VDD.n535 VSS 0.0147f
C1395 VDD.t95 VSS 0.01535f
C1396 VDD.n536 VSS 0.02464f
C1397 VDD.n537 VSS 0.0147f
C1398 VDD.n539 VSS 0.02306f
C1399 VDD.n540 VSS 0.03911f
C1400 VDD.t93 VSS 0.09216f
C1401 VDD.n541 VSS 0.02588f
C1402 VDD.n542 VSS 0.0147f
C1403 VDD.n543 VSS 0.0147f
C1404 VDD.n544 VSS 0.02588f
C1405 VDD.t58 VSS 0.09216f
C1406 VDD.n545 VSS 0.02588f
C1407 VDD.n546 VSS 0.0147f
C1408 VDD.n547 VSS 0.0147f
C1409 VDD.n548 VSS 0.02588f
C1410 VDD.t46 VSS 0.09216f
C1411 VDD.n549 VSS 0.02588f
C1412 VDD.n550 VSS 0.0147f
C1413 VDD.n551 VSS 0.0147f
C1414 VDD.n552 VSS 0.02588f
C1415 VDD.t84 VSS 0.09216f
C1416 VDD.n553 VSS 0.02588f
C1417 VDD.n554 VSS 0.01526f
C1418 VDD.n559 VSS 0.2614f
C1419 VDD.t47 VSS 0.09455f
C1420 VDD.n621 VSS 0.1891f
C1421 VDD.t8 VSS 0.09455f
C1422 VDD.n628 VSS 0.1891f
C1423 VDD.t0 VSS 0.09455f
C1424 VDD.n635 VSS 0.1891f
C1425 VDD.t30 VSS 0.09455f
C1426 VDD.n642 VSS 0.18771f
C1427 VDD.n646 VSS 0.1891f
C1428 VDD.t11 VSS 0.09455f
C1429 VDD.n650 VSS 0.16824f
C1430 VDD.n654 VSS 0.1891f
C1431 VDD.t44 VSS 0.09455f
C1432 VDD.n658 VSS 0.27531f
C1433 VDD.n721 VSS 0.22247f
C1434 VDD.n727 VSS 0.11541f
C1435 VDD.n733 VSS 0.1891f
C1436 VDD.n739 VSS 0.09594f
C1437 VDD.n745 VSS 0.17102f
C1438 VDD.n746 VSS 0.1891f
C1439 VDD.n752 VSS 0.11263f
C1440 VDD.n758 VSS 0.15156f
C1441 VDD.n759 VSS 0.1891f
C1442 VDD.n765 VSS 0.13209f
C1443 VDD.n771 VSS 0.13209f
C1444 VDD.n772 VSS 0.1891f
C1445 VDD.n778 VSS 0.15156f
C1446 VDD.n784 VSS 0.11263f
C1447 VDD.n785 VSS 0.1891f
C1448 VDD.n791 VSS 0.17102f
C1449 VDD.n798 VSS 0.31424f
C1450 VDD.n802 VSS 0.0185f
C1451 VDD.n803 VSS 0.02626f
C1452 VDD.n804 VSS 0.2902f
C1453 VDD.n805 VSS 0.2911f
C1454 VDD.n806 VSS 0.03622f
C1455 VDD.n807 VSS 0.05112f
C1456 VDD.n808 VSS 0.03362f
C1457 VDD.n809 VSS 0.13834f
C1458 a_8862_4192.t3 VSS 0.01275f
C1459 a_8862_4192.t16 VSS 0.01275f
C1460 a_8862_4192.t15 VSS 0.01275f
C1461 a_8862_4192.n0 VSS 0.03008f
C1462 a_8862_4192.t8 VSS 0.01275f
C1463 a_8862_4192.t7 VSS 0.01275f
C1464 a_8862_4192.n1 VSS 0.02863f
C1465 a_8862_4192.n2 VSS 0.20152f
C1466 a_8862_4192.t4 VSS 0.01275f
C1467 a_8862_4192.t27 VSS 0.01275f
C1468 a_8862_4192.n3 VSS 0.02863f
C1469 a_8862_4192.n4 VSS 0.11251f
C1470 a_8862_4192.t2 VSS 0.01275f
C1471 a_8862_4192.t1 VSS 0.01275f
C1472 a_8862_4192.n5 VSS 0.02863f
C1473 a_8862_4192.n6 VSS 0.11251f
C1474 a_8862_4192.t6 VSS 0.01275f
C1475 a_8862_4192.t5 VSS 0.01275f
C1476 a_8862_4192.n7 VSS 0.02863f
C1477 a_8862_4192.n8 VSS 0.11251f
C1478 a_8862_4192.t20 VSS 0.01275f
C1479 a_8862_4192.t18 VSS 0.01275f
C1480 a_8862_4192.n9 VSS 0.02863f
C1481 a_8862_4192.n10 VSS 0.11251f
C1482 a_8862_4192.t12 VSS 0.01275f
C1483 a_8862_4192.t10 VSS 0.01275f
C1484 a_8862_4192.n11 VSS 0.02863f
C1485 a_8862_4192.n12 VSS 0.21808f
C1486 a_8862_4192.t22 VSS 0.01275f
C1487 a_8862_4192.t21 VSS 0.01275f
C1488 a_8862_4192.n13 VSS 0.02863f
C1489 a_8862_4192.n14 VSS 0.21808f
C1490 a_8862_4192.t26 VSS 0.01275f
C1491 a_8862_4192.t25 VSS 0.01275f
C1492 a_8862_4192.n15 VSS 0.02863f
C1493 a_8862_4192.n16 VSS 0.11251f
C1494 a_8862_4192.t14 VSS 0.01275f
C1495 a_8862_4192.t13 VSS 0.01275f
C1496 a_8862_4192.n17 VSS 0.02863f
C1497 a_8862_4192.n18 VSS 0.11251f
C1498 a_8862_4192.t24 VSS 0.01275f
C1499 a_8862_4192.t23 VSS 0.01275f
C1500 a_8862_4192.n19 VSS 0.03008f
C1501 a_8862_4192.t19 VSS 0.01275f
C1502 a_8862_4192.t17 VSS 0.01275f
C1503 a_8862_4192.n20 VSS 0.02863f
C1504 a_8862_4192.n21 VSS 0.20152f
C1505 a_8862_4192.t11 VSS 0.01275f
C1506 a_8862_4192.t9 VSS 0.01275f
C1507 a_8862_4192.n22 VSS 0.02863f
C1508 a_8862_4192.n23 VSS 0.11251f
C1509 a_8862_4192.n24 VSS 0.11251f
C1510 a_8862_4192.n25 VSS 0.02863f
C1511 a_8862_4192.t0 VSS 0.01275f
C1512 EN.t47 VSS 0.24131f
C1513 EN.t50 VSS 0.24011f
C1514 EN.n0 VSS 0.47355f
C1515 EN.t17 VSS 0.24011f
C1516 EN.n1 VSS 0.24683f
C1517 EN.t19 VSS 0.24011f
C1518 EN.n2 VSS 0.42772f
C1519 EN.t69 VSS 0.24131f
C1520 EN.t71 VSS 0.24011f
C1521 EN.n3 VSS 0.47355f
C1522 EN.t44 VSS 0.24011f
C1523 EN.n4 VSS 0.24683f
C1524 EN.t46 VSS 0.24011f
C1525 EN.n5 VSS 0.40435f
C1526 EN.n6 VSS 0.39676f
C1527 EN.t91 VSS 0.24131f
C1528 EN.t0 VSS 0.24011f
C1529 EN.n7 VSS 0.47355f
C1530 EN.t61 VSS 0.24011f
C1531 EN.n8 VSS 0.24683f
C1532 EN.t65 VSS 0.24011f
C1533 EN.n9 VSS 0.40435f
C1534 EN.n10 VSS 0.40266f
C1535 EN.t85 VSS 0.24131f
C1536 EN.t87 VSS 0.24011f
C1537 EN.n11 VSS 0.47355f
C1538 EN.t56 VSS 0.24011f
C1539 EN.n12 VSS 0.24683f
C1540 EN.t57 VSS 0.24011f
C1541 EN.n13 VSS 0.40435f
C1542 EN.n14 VSS 0.40266f
C1543 EN.t41 VSS 0.24131f
C1544 EN.t45 VSS 0.24011f
C1545 EN.n15 VSS 0.47355f
C1546 EN.t9 VSS 0.24011f
C1547 EN.n16 VSS 0.24683f
C1548 EN.t10 VSS 0.24011f
C1549 EN.n17 VSS 0.40435f
C1550 EN.n18 VSS 0.28088f
C1551 EN.t66 VSS 0.24147f
C1552 EN.t21 VSS 0.24024f
C1553 EN.n19 VSS 0.58221f
C1554 EN.t13 VSS 0.24024f
C1555 EN.n20 VSS 0.34898f
C1556 EN.t48 VSS 0.24024f
C1557 EN.n21 VSS 0.57396f
C1558 EN.t72 VSS 0.24248f
C1559 EN.t70 VSS 0.24024f
C1560 EN.n22 VSS 0.77242f
C1561 EN.t22 VSS 0.24024f
C1562 EN.n23 VSS 0.34898f
C1563 EN.t20 VSS 0.24024f
C1564 EN.n24 VSS 0.41089f
C1565 EN.n25 VSS 0.59874f
C1566 EN.t35 VSS 0.24147f
C1567 EN.t90 VSS 0.24024f
C1568 EN.n26 VSS 0.58221f
C1569 EN.t78 VSS 0.24024f
C1570 EN.n27 VSS 0.34898f
C1571 EN.t16 VSS 0.24024f
C1572 EN.n28 VSS 0.50657f
C1573 EN.n29 VSS 0.42968f
C1574 EN.t39 VSS 0.24248f
C1575 EN.t37 VSS 0.24024f
C1576 EN.n30 VSS 0.77242f
C1577 EN.t86 VSS 0.24024f
C1578 EN.n31 VSS 0.34898f
C1579 EN.t81 VSS 0.24024f
C1580 EN.n32 VSS 0.41089f
C1581 EN.n33 VSS 0.33415f
C1582 EN.t34 VSS 0.24147f
C1583 EN.t89 VSS 0.24024f
C1584 EN.n34 VSS 0.58221f
C1585 EN.t77 VSS 0.24024f
C1586 EN.n35 VSS 0.34898f
C1587 EN.t15 VSS 0.24024f
C1588 EN.n36 VSS 0.50657f
C1589 EN.n37 VSS 0.42836f
C1590 EN.t38 VSS 0.24248f
C1591 EN.t33 VSS 0.24024f
C1592 EN.n38 VSS 0.77242f
C1593 EN.t84 VSS 0.24024f
C1594 EN.n39 VSS 0.34898f
C1595 EN.t76 VSS 0.24024f
C1596 EN.n40 VSS 0.36635f
C1597 EN.t83 VSS 0.24248f
C1598 EN.t60 VSS 0.24024f
C1599 EN.n41 VSS 0.77242f
C1600 EN.t64 VSS 0.24024f
C1601 EN.n42 VSS 0.34898f
C1602 EN.t51 VSS 0.24024f
C1603 EN.n43 VSS 0.62852f
C1604 EN.t25 VSS 0.24147f
C1605 EN.t27 VSS 0.24024f
C1606 EN.n44 VSS 0.58221f
C1607 EN.t30 VSS 0.24024f
C1608 EN.n45 VSS 0.34898f
C1609 EN.t8 VSS 0.24024f
C1610 EN.n46 VSS 0.34898f
C1611 EN.t68 VSS 0.24024f
C1612 EN.n47 VSS 0.34898f
C1613 EN.t43 VSS 0.24024f
C1614 EN.n48 VSS 0.46467f
C1615 EN.n49 VSS 0.70337f
C1616 EN.t82 VSS 0.24248f
C1617 EN.t59 VSS 0.24024f
C1618 EN.n50 VSS 0.77242f
C1619 EN.t62 VSS 0.24024f
C1620 EN.n51 VSS 0.34898f
C1621 EN.t49 VSS 0.24024f
C1622 EN.n52 VSS 0.34898f
C1623 EN.t14 VSS 0.24024f
C1624 EN.n53 VSS 0.34898f
C1625 EN.t12 VSS 0.24024f
C1626 EN.n54 VSS 0.36895f
C1627 EN.n55 VSS 0.29233f
C1628 EN.t24 VSS 0.24147f
C1629 EN.t26 VSS 0.24024f
C1630 EN.n56 VSS 0.58221f
C1631 EN.t29 VSS 0.24024f
C1632 EN.n57 VSS 0.34898f
C1633 EN.t7 VSS 0.24024f
C1634 EN.n58 VSS 0.34898f
C1635 EN.t67 VSS 0.24024f
C1636 EN.n59 VSS 0.34898f
C1637 EN.t42 VSS 0.24024f
C1638 EN.n60 VSS 0.46467f
C1639 EN.n61 VSS 0.38783f
C1640 EN.t55 VSS 0.24248f
C1641 EN.t28 VSS 0.24024f
C1642 EN.n62 VSS 0.77242f
C1643 EN.t32 VSS 0.24024f
C1644 EN.n63 VSS 0.34898f
C1645 EN.t18 VSS 0.24024f
C1646 EN.n64 VSS 0.34898f
C1647 EN.t80 VSS 0.24024f
C1648 EN.n65 VSS 0.34898f
C1649 EN.t75 VSS 0.24024f
C1650 EN.n66 VSS 0.36895f
C1651 EN.n67 VSS 0.29233f
C1652 EN.t1 VSS 0.24147f
C1653 EN.t2 VSS 0.24024f
C1654 EN.n68 VSS 0.58221f
C1655 EN.t3 VSS 0.24024f
C1656 EN.n69 VSS 0.34898f
C1657 EN.t74 VSS 0.24024f
C1658 EN.n70 VSS 0.34898f
C1659 EN.t40 VSS 0.24024f
C1660 EN.n71 VSS 0.34898f
C1661 EN.t6 VSS 0.24024f
C1662 EN.n72 VSS 0.46467f
C1663 EN.n73 VSS 0.38783f
C1664 EN.t23 VSS 0.24248f
C1665 EN.t4 VSS 0.24024f
C1666 EN.n74 VSS 0.77242f
C1667 EN.t5 VSS 0.24024f
C1668 EN.n75 VSS 0.34898f
C1669 EN.t88 VSS 0.24024f
C1670 EN.n76 VSS 0.34898f
C1671 EN.t54 VSS 0.24024f
C1672 EN.n77 VSS 0.34898f
C1673 EN.t52 VSS 0.24024f
C1674 EN.n78 VSS 0.36895f
C1675 EN.n79 VSS 0.29233f
C1676 EN.t73 VSS 0.24348f
C1677 EN.t53 VSS 0.24024f
C1678 EN.n80 VSS 0.96263f
C1679 EN.t11 VSS 0.24024f
C1680 EN.n81 VSS 0.34898f
C1681 EN.t79 VSS 0.24024f
C1682 EN.n82 VSS 0.46467f
C1683 EN.n83 VSS 1.61336f
C1684 EN.n84 VSS 1.57146f
C1685 EN.n85 VSS 0.24599f
C1686 EN.n86 VSS 0.23361f
C1687 EN.t58 VSS 0.24131f
C1688 EN.t63 VSS 0.24011f
C1689 EN.n87 VSS 0.47355f
C1690 EN.t31 VSS 0.24011f
C1691 EN.n88 VSS 0.24683f
C1692 EN.t36 VSS 0.24011f
C1693 EN.n89 VSS 0.37076f
C1694 EN.n90 VSS 1.23156f
.ends

