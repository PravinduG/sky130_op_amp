magic
tech sky130A
magscale 1 2
timestamp 1761058420
<< pwell >>
rect -297 1586 297 1672
rect -297 -1586 -211 1586
rect 211 -1586 297 1586
rect -297 -1672 297 -1586
<< psubdiff >>
rect -271 1612 -153 1646
rect -119 1612 -85 1646
rect -51 1612 -17 1646
rect 17 1612 51 1646
rect 85 1612 119 1646
rect 153 1612 271 1646
rect -271 1547 -237 1612
rect 237 1547 271 1612
rect -271 1479 -237 1513
rect -271 1411 -237 1445
rect -271 1343 -237 1377
rect -271 1275 -237 1309
rect -271 1207 -237 1241
rect -271 1139 -237 1173
rect -271 1071 -237 1105
rect -271 1003 -237 1037
rect -271 935 -237 969
rect -271 867 -237 901
rect -271 799 -237 833
rect -271 731 -237 765
rect -271 663 -237 697
rect -271 595 -237 629
rect -271 527 -237 561
rect -271 459 -237 493
rect -271 391 -237 425
rect -271 323 -237 357
rect -271 255 -237 289
rect -271 187 -237 221
rect -271 119 -237 153
rect -271 51 -237 85
rect -271 -17 -237 17
rect -271 -85 -237 -51
rect -271 -153 -237 -119
rect -271 -221 -237 -187
rect -271 -289 -237 -255
rect -271 -357 -237 -323
rect -271 -425 -237 -391
rect -271 -493 -237 -459
rect -271 -561 -237 -527
rect -271 -629 -237 -595
rect -271 -697 -237 -663
rect -271 -765 -237 -731
rect -271 -833 -237 -799
rect -271 -901 -237 -867
rect -271 -969 -237 -935
rect -271 -1037 -237 -1003
rect -271 -1105 -237 -1071
rect -271 -1173 -237 -1139
rect -271 -1241 -237 -1207
rect -271 -1309 -237 -1275
rect -271 -1377 -237 -1343
rect -271 -1445 -237 -1411
rect -271 -1513 -237 -1479
rect 237 1479 271 1513
rect 237 1411 271 1445
rect 237 1343 271 1377
rect 237 1275 271 1309
rect 237 1207 271 1241
rect 237 1139 271 1173
rect 237 1071 271 1105
rect 237 1003 271 1037
rect 237 935 271 969
rect 237 867 271 901
rect 237 799 271 833
rect 237 731 271 765
rect 237 663 271 697
rect 237 595 271 629
rect 237 527 271 561
rect 237 459 271 493
rect 237 391 271 425
rect 237 323 271 357
rect 237 255 271 289
rect 237 187 271 221
rect 237 119 271 153
rect 237 51 271 85
rect 237 -17 271 17
rect 237 -85 271 -51
rect 237 -153 271 -119
rect 237 -221 271 -187
rect 237 -289 271 -255
rect 237 -357 271 -323
rect 237 -425 271 -391
rect 237 -493 271 -459
rect 237 -561 271 -527
rect 237 -629 271 -595
rect 237 -697 271 -663
rect 237 -765 271 -731
rect 237 -833 271 -799
rect 237 -901 271 -867
rect 237 -969 271 -935
rect 237 -1037 271 -1003
rect 237 -1105 271 -1071
rect 237 -1173 271 -1139
rect 237 -1241 271 -1207
rect 237 -1309 271 -1275
rect 237 -1377 271 -1343
rect 237 -1445 271 -1411
rect 237 -1513 271 -1479
rect -271 -1612 -237 -1547
rect 237 -1612 271 -1547
rect -271 -1646 -153 -1612
rect -119 -1646 -85 -1612
rect -51 -1646 -17 -1612
rect 17 -1646 51 -1612
rect 85 -1646 119 -1612
rect 153 -1646 271 -1612
<< psubdiffcont >>
rect -153 1612 -119 1646
rect -85 1612 -51 1646
rect -17 1612 17 1646
rect 51 1612 85 1646
rect 119 1612 153 1646
rect -271 1513 -237 1547
rect -271 1445 -237 1479
rect -271 1377 -237 1411
rect -271 1309 -237 1343
rect -271 1241 -237 1275
rect -271 1173 -237 1207
rect -271 1105 -237 1139
rect -271 1037 -237 1071
rect -271 969 -237 1003
rect -271 901 -237 935
rect -271 833 -237 867
rect -271 765 -237 799
rect -271 697 -237 731
rect -271 629 -237 663
rect -271 561 -237 595
rect -271 493 -237 527
rect -271 425 -237 459
rect -271 357 -237 391
rect -271 289 -237 323
rect -271 221 -237 255
rect -271 153 -237 187
rect -271 85 -237 119
rect -271 17 -237 51
rect -271 -51 -237 -17
rect -271 -119 -237 -85
rect -271 -187 -237 -153
rect -271 -255 -237 -221
rect -271 -323 -237 -289
rect -271 -391 -237 -357
rect -271 -459 -237 -425
rect -271 -527 -237 -493
rect -271 -595 -237 -561
rect -271 -663 -237 -629
rect -271 -731 -237 -697
rect -271 -799 -237 -765
rect -271 -867 -237 -833
rect -271 -935 -237 -901
rect -271 -1003 -237 -969
rect -271 -1071 -237 -1037
rect -271 -1139 -237 -1105
rect -271 -1207 -237 -1173
rect -271 -1275 -237 -1241
rect -271 -1343 -237 -1309
rect -271 -1411 -237 -1377
rect -271 -1479 -237 -1445
rect -271 -1547 -237 -1513
rect 237 1513 271 1547
rect 237 1445 271 1479
rect 237 1377 271 1411
rect 237 1309 271 1343
rect 237 1241 271 1275
rect 237 1173 271 1207
rect 237 1105 271 1139
rect 237 1037 271 1071
rect 237 969 271 1003
rect 237 901 271 935
rect 237 833 271 867
rect 237 765 271 799
rect 237 697 271 731
rect 237 629 271 663
rect 237 561 271 595
rect 237 493 271 527
rect 237 425 271 459
rect 237 357 271 391
rect 237 289 271 323
rect 237 221 271 255
rect 237 153 271 187
rect 237 85 271 119
rect 237 17 271 51
rect 237 -51 271 -17
rect 237 -119 271 -85
rect 237 -187 271 -153
rect 237 -255 271 -221
rect 237 -323 271 -289
rect 237 -391 271 -357
rect 237 -459 271 -425
rect 237 -527 271 -493
rect 237 -595 271 -561
rect 237 -663 271 -629
rect 237 -731 271 -697
rect 237 -799 271 -765
rect 237 -867 271 -833
rect 237 -935 271 -901
rect 237 -1003 271 -969
rect 237 -1071 271 -1037
rect 237 -1139 271 -1105
rect 237 -1207 271 -1173
rect 237 -1275 271 -1241
rect 237 -1343 271 -1309
rect 237 -1411 271 -1377
rect 237 -1479 271 -1445
rect 237 -1547 271 -1513
rect -153 -1646 -119 -1612
rect -85 -1646 -51 -1612
rect -17 -1646 17 -1612
rect 51 -1646 85 -1612
rect 119 -1646 153 -1612
<< xpolycontact >>
rect -141 1084 141 1516
rect -141 -1516 141 -1084
<< xpolyres >>
rect -141 -1084 141 1084
<< locali >>
rect -271 1612 -153 1646
rect -119 1612 -85 1646
rect -51 1612 -17 1646
rect 17 1612 51 1646
rect 85 1612 119 1646
rect 153 1612 271 1646
rect -271 1547 -237 1612
rect 237 1547 271 1612
rect -271 1479 -237 1513
rect -271 1411 -237 1445
rect -271 1343 -237 1377
rect -271 1275 -237 1309
rect -271 1207 -237 1241
rect -271 1139 -237 1173
rect -271 1071 -237 1105
rect 237 1479 271 1513
rect 237 1411 271 1445
rect 237 1343 271 1377
rect 237 1275 271 1309
rect 237 1207 271 1241
rect 237 1139 271 1173
rect -271 1003 -237 1037
rect -271 935 -237 969
rect -271 867 -237 901
rect -271 799 -237 833
rect -271 731 -237 765
rect -271 663 -237 697
rect -271 595 -237 629
rect -271 527 -237 561
rect -271 459 -237 493
rect -271 391 -237 425
rect -271 323 -237 357
rect -271 255 -237 289
rect -271 187 -237 221
rect -271 119 -237 153
rect -271 51 -237 85
rect -271 -17 -237 17
rect -271 -85 -237 -51
rect -271 -153 -237 -119
rect -271 -221 -237 -187
rect -271 -289 -237 -255
rect -271 -357 -237 -323
rect -271 -425 -237 -391
rect -271 -493 -237 -459
rect -271 -561 -237 -527
rect -271 -629 -237 -595
rect -271 -697 -237 -663
rect -271 -765 -237 -731
rect -271 -833 -237 -799
rect -271 -901 -237 -867
rect -271 -969 -237 -935
rect -271 -1037 -237 -1003
rect -271 -1105 -237 -1071
rect 237 1071 271 1105
rect 237 1003 271 1037
rect 237 935 271 969
rect 237 867 271 901
rect 237 799 271 833
rect 237 731 271 765
rect 237 663 271 697
rect 237 595 271 629
rect 237 527 271 561
rect 237 459 271 493
rect 237 391 271 425
rect 237 323 271 357
rect 237 255 271 289
rect 237 187 271 221
rect 237 119 271 153
rect 237 51 271 85
rect 237 -17 271 17
rect 237 -85 271 -51
rect 237 -153 271 -119
rect 237 -221 271 -187
rect 237 -289 271 -255
rect 237 -357 271 -323
rect 237 -425 271 -391
rect 237 -493 271 -459
rect 237 -561 271 -527
rect 237 -629 271 -595
rect 237 -697 271 -663
rect 237 -765 271 -731
rect 237 -833 271 -799
rect 237 -901 271 -867
rect 237 -969 271 -935
rect 237 -1037 271 -1003
rect -271 -1173 -237 -1139
rect -271 -1241 -237 -1207
rect -271 -1309 -237 -1275
rect -271 -1377 -237 -1343
rect -271 -1445 -237 -1411
rect -271 -1513 -237 -1479
rect 237 -1105 271 -1071
rect 237 -1173 271 -1139
rect 237 -1241 271 -1207
rect 237 -1309 271 -1275
rect 237 -1377 271 -1343
rect 237 -1445 271 -1411
rect 237 -1513 271 -1479
rect -271 -1612 -237 -1547
rect 237 -1612 271 -1547
rect -271 -1646 -153 -1612
rect -119 -1646 -85 -1612
rect -51 -1646 -17 -1612
rect 17 -1646 51 -1612
rect 85 -1646 119 -1612
rect 153 -1646 271 -1612
<< viali >>
rect -125 1102 125 1496
rect -125 -1497 125 -1103
<< metal1 >>
rect -131 1496 131 1510
rect -131 1102 -125 1496
rect 125 1102 131 1496
rect -131 1089 131 1102
rect -131 -1103 131 -1089
rect -131 -1497 -125 -1103
rect 125 -1497 131 -1103
rect -131 -1510 131 -1497
<< properties >>
string FIXED_BBOX -254 -1629 254 1629
<< end >>
