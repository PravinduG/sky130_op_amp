** sch_path: /foss/designs/sky130_op_amp/runs/RUN_2025-10-21_18-07-48/parameters/offset_params/run_05/sky130_op_amp_tb.sch
**.subckt sky130_op_amp_tb
C1 Vout VSS 2.5e-11 m=1
Vdm net2 GND ac 1
Vcm net1 GND 0.9
I0 VDD IBIAS 4.9999999999999996e-06
E2 VN net1 net2 GND -0.5
E1 VP net1 net2 GND 0.5
V0 VSS GND 0
V4 VDD GND CACE{vdd}
x1 VDD IBIAS VN VP Vout VDD VSS sky130_op_amp
**** begin user architecture code


.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt

.include /foss/designs/sky130_op_amp/netlist/rcx/sky130_op_amp.spice

.temp 27

.option SEED=12345

* Flag unsafe operating conditions (exceeds models' specified limits)
.option warn=1




.control
*---------------------------------------
* AC Analysis (DC gain, UGF, Phase Margin)
*---------------------------------------
ac dec 20 1k 100e6
let vout_mag = abs(v(Vout))
let vout_phase = phase(v(Vout))*180/pi
meas ac a0 find vout_mag at=1k
meas ac ugf when vout_mag=1 fall=1
meas ac pm find 180+vout_phase when vout_mag=1

*---------------------------------------
* Output Offset (Vin = 0.9V)
*---------------------------------------
dc Vcm 0.9 0.9 0.1
meas dc vout_offset find v(Vout) at=0.9

*---------------------------------------
* Input Offset (Vout = 0.9V)
*---------------------------------------
dc Vcm 0.85 0.95 0.001
meas dc vin_offset when v(Vout)=0.9

*---------------------------------------
* Slew Rate (Transient)
*---------------------------------------
Vstep VIN GND PULSE(0.9 1.1 1u 0.1u 0.1u 4u 8u)
tran 0.05u 10u
meas tran sr_pos max deriv(v(Vout))

alter Vstep PULSE(0.9 0.7 1u 0.1u 0.1u 4u 8u)
tran 0.05u 10u
meas tran sr_neg min deriv(v(Vout))

*---------------------------------------
* Supply Current (Enabled/Disabled)
*---------------------------------------
dc Ven 1.8 1.8 0.1
meas dc idd_enabled find -i(Vdd)

alter Ven 0
dc Ven 0 0 0.1
meas dc idd_disabled find -i(Vdd)

*---------------------------------------
* Echo all measurements
*---------------------------------------
echo $&a0 $&ugf $&pm $&vout_offset $&vin_offset $&sr_pos $&sr_neg $&idd_enabled $&idd_disabled > /foss/designs/sky130_op_amp/runs/RUN_2025-10-21_18-07-48/parameters/offset_params/run_05/sky130_op_amp_tb_5.data
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
